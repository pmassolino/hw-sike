----------------------------------------------------------------------------------
-- Implementation by Pedro Maat C. Massolino,
-- hereby denoted as "the implementer".
--
-- To the extent possible under law, the implementer has waived all copyright
-- and related or neighboring rights to the source code in this file.
-- http://creativecommons.org/publicdomain/zero/1.0/
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity carmela_state_machine_v128 is
    Port (
        clk : in std_logic;
        rstn : in std_logic;
        instruction_values_valid : in std_logic;
        instruction_type : in std_logic_vector(3 downto 0);
        operands_size : in std_logic_vector(2 downto 0);
        prime_line_equal_one : in std_logic_vector(1 downto 0);
        penultimate_operation : in std_logic;
        sm_rotation_size : out std_logic_vector(1 downto 0);
        sm_circular_shift_enable : out std_logic;
        sel_address_a : out std_logic;
        sel_address_b_prime : out std_logic_vector(1 downto 0);
        sm_specific_mac_address_a : out std_logic_vector(2 downto 0);
        sm_specific_mac_address_b : out std_logic_vector(2 downto 0);
        sm_specific_mac_address_o : out std_logic_vector(2 downto 0);
        sm_specific_mac_next_address_o : out std_logic_vector(2 downto 0);
        mac_enable_signed_a : out std_logic;
        mac_enable_signed_b : out std_logic;
        mac_sel_load_reg_a : out std_logic_vector(1 downto 0);
        mac_clear_reg_b : out std_logic;
        mac_clear_reg_acc : out std_logic;
        mac_sel_shift_reg_o : out std_logic;
        mac_enable_update_reg_s : out std_logic;
        mac_sel_reg_s_reg_o_sign : out std_logic;
        mac_reg_s_reg_o_positive : out std_logic;
        sm_sign_a_mode : out std_logic;
        sm_mac_operation_mode : out std_logic_vector(1 downto 0);
        mac_enable_reg_s_mask : out std_logic;
        mac_subtraction_reg_a_b : out std_logic;
        mac_sel_multiply_two_a_b : out std_logic;
        mac_sel_reg_y_output : out std_logic;
        sm_mac_write_enable_output : out std_logic;
        mac_memory_double_mode : out std_logic;
        mac_memory_only_write_mode : out std_logic;
        base_address_generator_o_increment_previous_address : out std_logic;
        sm_free_flag : out std_logic
    );
end carmela_state_machine_v128;

architecture behavioral of carmela_state_machine_v128 is

type state is (reset, decode_instruction,
-- 0000 multiplication with no reduction
multiplication_direct_0,
multiplication_direct_2, multiplication_direct_3, multiplication_direct_4, multiplication_direct_5,
multiplication_direct_7, multiplication_direct_8, multiplication_direct_9, multiplication_direct_10, multiplication_direct_11, multiplication_direct_12, multiplication_direct_13, multiplication_direct_14,
multiplication_direct_16, multiplication_direct_17, multiplication_direct_18, multiplication_direct_19, multiplication_direct_20, multiplication_direct_21, multiplication_direct_22, multiplication_direct_23, multiplication_direct_24, multiplication_direct_25, multiplication_direct_26, multiplication_direct_27,
multiplication_direct_29, multiplication_direct_30, multiplication_direct_31, multiplication_direct_32, multiplication_direct_33, multiplication_direct_34, multiplication_direct_35, multiplication_direct_36, multiplication_direct_37, multiplication_direct_38, multiplication_direct_39, multiplication_direct_40, multiplication_direct_41, multiplication_direct_42, multiplication_direct_43, multiplication_direct_44, multiplication_direct_45,
multiplication_direct_47, multiplication_direct_48, multiplication_direct_49, multiplication_direct_50, multiplication_direct_51, multiplication_direct_52, multiplication_direct_53, multiplication_direct_54, multiplication_direct_55, multiplication_direct_56, multiplication_direct_57, multiplication_direct_58, multiplication_direct_59, multiplication_direct_60, multiplication_direct_61, multiplication_direct_62, multiplication_direct_63, multiplication_direct_64, multiplication_direct_65, multiplication_direct_66, multiplication_direct_67, multiplication_direct_68, multiplication_direct_69,
multiplication_direct_71, multiplication_direct_72, multiplication_direct_73, multiplication_direct_74, multiplication_direct_75, multiplication_direct_76, multiplication_direct_77, multiplication_direct_78, multiplication_direct_79, multiplication_direct_80, multiplication_direct_81, multiplication_direct_82, multiplication_direct_83, multiplication_direct_84, multiplication_direct_85, multiplication_direct_86, multiplication_direct_87, multiplication_direct_88, multiplication_direct_89, multiplication_direct_90, multiplication_direct_91, multiplication_direct_92, multiplication_direct_93, multiplication_direct_94, multiplication_direct_95, multiplication_direct_96, multiplication_direct_97, multiplication_direct_98, multiplication_direct_99, multiplication_direct_100,
multiplication_direct_102, multiplication_direct_103, multiplication_direct_104, multiplication_direct_105, multiplication_direct_106, multiplication_direct_107, multiplication_direct_108, multiplication_direct_109, multiplication_direct_110, multiplication_direct_111, multiplication_direct_112, multiplication_direct_113, multiplication_direct_114, multiplication_direct_115, multiplication_direct_116, multiplication_direct_117, multiplication_direct_118, multiplication_direct_119, multiplication_direct_120, multiplication_direct_121, multiplication_direct_122, multiplication_direct_123, multiplication_direct_124, multiplication_direct_125, multiplication_direct_126, multiplication_direct_127, multiplication_direct_128, multiplication_direct_129, multiplication_direct_130, multiplication_direct_131, multiplication_direct_132, multiplication_direct_133, multiplication_direct_134, multiplication_direct_135, multiplication_direct_136, multiplication_direct_137, multiplication_direct_138, multiplication_direct_139,
-- 0001 square with no reduction
square_direct_0,
square_direct_2, square_direct_3, square_direct_4,
square_direct_6, square_direct_7, square_direct_8, square_direct_9, square_direct_10,
square_direct_12, square_direct_13, square_direct_14, square_direct_15, square_direct_16, square_direct_17, square_direct_18,
square_direct_20, square_direct_21, square_direct_22, square_direct_23, square_direct_24, square_direct_25, square_direct_26, square_direct_27, square_direct_28, square_direct_29,
square_direct_31, square_direct_32, square_direct_33, square_direct_34, square_direct_35, square_direct_36, square_direct_37, square_direct_38, square_direct_39, square_direct_40, square_direct_41, square_direct_42, square_direct_43,
square_direct_45, square_direct_46, square_direct_47, square_direct_48, square_direct_49, square_direct_50, square_direct_51, square_direct_52, square_direct_53, square_direct_54, square_direct_55, square_direct_56, square_direct_57, square_direct_58, square_direct_59, square_direct_60, square_direct_61,
square_direct_63, square_direct_64, square_direct_65, square_direct_66, square_direct_67, square_direct_68, square_direct_69, square_direct_70, square_direct_71, square_direct_72, square_direct_73, square_direct_74, square_direct_75, square_direct_76, square_direct_77, square_direct_78, square_direct_79, square_direct_80, square_direct_81, square_direct_82, square_direct_83,
-- 0010 multiplication with reduction and prime line not equal to 1
multiplication_with_reduction_0, multiplication_with_reduction_1, multiplication_with_reduction_2, multiplication_with_reduction_3,
multiplication_with_reduction_5, multiplication_with_reduction_6, multiplication_with_reduction_7, multiplication_with_reduction_8, multiplication_with_reduction_9, multiplication_with_reduction_10, multiplication_with_reduction_11, multiplication_with_reduction_12, multiplication_with_reduction_13, multiplication_with_reduction_14,
multiplication_with_reduction_16, multiplication_with_reduction_17, multiplication_with_reduction_18, multiplication_with_reduction_19, multiplication_with_reduction_20, multiplication_with_reduction_21, multiplication_with_reduction_22, multiplication_with_reduction_23, multiplication_with_reduction_24, multiplication_with_reduction_25, multiplication_with_reduction_26, multiplication_with_reduction_27, multiplication_with_reduction_28, multiplication_with_reduction_29, multiplication_with_reduction_30, multiplication_with_reduction_31, multiplication_with_reduction_32,
multiplication_with_reduction_34, multiplication_with_reduction_35, multiplication_with_reduction_36, multiplication_with_reduction_37, multiplication_with_reduction_38, multiplication_with_reduction_39, multiplication_with_reduction_40, multiplication_with_reduction_41, multiplication_with_reduction_42, multiplication_with_reduction_43, multiplication_with_reduction_44, multiplication_with_reduction_45, multiplication_with_reduction_46, multiplication_with_reduction_47, multiplication_with_reduction_48, multiplication_with_reduction_49, multiplication_with_reduction_50, multiplication_with_reduction_51, multiplication_with_reduction_52, multiplication_with_reduction_53, multiplication_with_reduction_54, multiplication_with_reduction_55, multiplication_with_reduction_56, multiplication_with_reduction_57, multiplication_with_reduction_58, 
multiplication_with_reduction_60, multiplication_with_reduction_61, multiplication_with_reduction_62, multiplication_with_reduction_63, multiplication_with_reduction_64,multiplication_with_reduction_65, multiplication_with_reduction_66, multiplication_with_reduction_67, multiplication_with_reduction_68, multiplication_with_reduction_69, multiplication_with_reduction_70, multiplication_with_reduction_71, multiplication_with_reduction_72, multiplication_with_reduction_73, multiplication_with_reduction_74,multiplication_with_reduction_75, multiplication_with_reduction_76, multiplication_with_reduction_77, multiplication_with_reduction_78, multiplication_with_reduction_79, multiplication_with_reduction_80, multiplication_with_reduction_81, multiplication_with_reduction_82, multiplication_with_reduction_83, multiplication_with_reduction_84, multiplication_with_reduction_85, multiplication_with_reduction_86, multiplication_with_reduction_87, multiplication_with_reduction_88, multiplication_with_reduction_89, multiplication_with_reduction_90, multiplication_with_reduction_91, multiplication_with_reduction_92, multiplication_with_reduction_93, multiplication_with_reduction_94, multiplication_with_reduction_96, multiplication_with_reduction_97, multiplication_with_reduction_98, multiplication_with_reduction_99, multiplication_with_reduction_100, multiplication_with_reduction_101, multiplication_with_reduction_102, multiplication_with_reduction_103, multiplication_with_reduction_104, multiplication_with_reduction_105, multiplication_with_reduction_106, multiplication_with_reduction_107, multiplication_with_reduction_108, multiplication_with_reduction_109, multiplication_with_reduction_110, multiplication_with_reduction_111, multiplication_with_reduction_112, multiplication_with_reduction_113, multiplication_with_reduction_114, multiplication_with_reduction_115, multiplication_with_reduction_116, multiplication_with_reduction_117, multiplication_with_reduction_118, multiplication_with_reduction_119, multiplication_with_reduction_120, multiplication_with_reduction_121, multiplication_with_reduction_122, multiplication_with_reduction_123, multiplication_with_reduction_124, multiplication_with_reduction_125, multiplication_with_reduction_126, multiplication_with_reduction_127, multiplication_with_reduction_128, multiplication_with_reduction_129, multiplication_with_reduction_130, multiplication_with_reduction_131, multiplication_with_reduction_132, multiplication_with_reduction_133, multiplication_with_reduction_134, multiplication_with_reduction_135, multiplication_with_reduction_136, multiplication_with_reduction_137, multiplication_with_reduction_138, multiplication_with_reduction_139, multiplication_with_reduction_140, multiplication_with_reduction_141, multiplication_with_reduction_142,
multiplication_with_reduction_144, multiplication_with_reduction_145, multiplication_with_reduction_146, multiplication_with_reduction_147, multiplication_with_reduction_148, multiplication_with_reduction_149, multiplication_with_reduction_150, multiplication_with_reduction_151, multiplication_with_reduction_152, multiplication_with_reduction_153, multiplication_with_reduction_154, multiplication_with_reduction_155, multiplication_with_reduction_156, multiplication_with_reduction_157, multiplication_with_reduction_158, multiplication_with_reduction_159, multiplication_with_reduction_160, multiplication_with_reduction_161, multiplication_with_reduction_162, multiplication_with_reduction_163, multiplication_with_reduction_164, multiplication_with_reduction_165, multiplication_with_reduction_166, multiplication_with_reduction_167, multiplication_with_reduction_168, multiplication_with_reduction_169, multiplication_with_reduction_170, multiplication_with_reduction_171, multiplication_with_reduction_172, multiplication_with_reduction_173, multiplication_with_reduction_174, multiplication_with_reduction_175, multiplication_with_reduction_176, multiplication_with_reduction_177, multiplication_with_reduction_178, multiplication_with_reduction_179, multiplication_with_reduction_180, multiplication_with_reduction_181, multiplication_with_reduction_182, multiplication_with_reduction_183, multiplication_with_reduction_184, multiplication_with_reduction_185, multiplication_with_reduction_186, multiplication_with_reduction_187, multiplication_with_reduction_188, multiplication_with_reduction_189, multiplication_with_reduction_190, multiplication_with_reduction_191, multiplication_with_reduction_192, multiplication_with_reduction_193, multiplication_with_reduction_194, multiplication_with_reduction_195, multiplication_with_reduction_196, multiplication_with_reduction_197, multiplication_with_reduction_198, multiplication_with_reduction_199, multiplication_with_reduction_200, multiplication_with_reduction_201, multiplication_with_reduction_202, multiplication_with_reduction_203, multiplication_with_reduction_204,
multiplication_with_reduction_206, multiplication_with_reduction_207, multiplication_with_reduction_208, multiplication_with_reduction_209, multiplication_with_reduction_210, multiplication_with_reduction_211, multiplication_with_reduction_212, multiplication_with_reduction_213, multiplication_with_reduction_214, multiplication_with_reduction_215, multiplication_with_reduction_216, multiplication_with_reduction_217, multiplication_with_reduction_218, multiplication_with_reduction_219, multiplication_with_reduction_220, multiplication_with_reduction_221, multiplication_with_reduction_222, multiplication_with_reduction_223, multiplication_with_reduction_224, multiplication_with_reduction_225, multiplication_with_reduction_226, multiplication_with_reduction_227, multiplication_with_reduction_228, multiplication_with_reduction_229, multiplication_with_reduction_230, multiplication_with_reduction_231, multiplication_with_reduction_232, multiplication_with_reduction_233, multiplication_with_reduction_234, multiplication_with_reduction_235, multiplication_with_reduction_236, multiplication_with_reduction_237, multiplication_with_reduction_238, multiplication_with_reduction_239, multiplication_with_reduction_240, multiplication_with_reduction_241, multiplication_with_reduction_242, multiplication_with_reduction_243, multiplication_with_reduction_244, multiplication_with_reduction_245, multiplication_with_reduction_246, multiplication_with_reduction_247, multiplication_with_reduction_248, multiplication_with_reduction_249, multiplication_with_reduction_250,multiplication_with_reduction_251, multiplication_with_reduction_252, multiplication_with_reduction_253, multiplication_with_reduction_254, multiplication_with_reduction_255, multiplication_with_reduction_256, multiplication_with_reduction_257, multiplication_with_reduction_258, multiplication_with_reduction_259, multiplication_with_reduction_260, multiplication_with_reduction_261, multiplication_with_reduction_262, multiplication_with_reduction_263, multiplication_with_reduction_264, multiplication_with_reduction_265, multiplication_with_reduction_266, multiplication_with_reduction_267, multiplication_with_reduction_268, multiplication_with_reduction_269, multiplication_with_reduction_270, multiplication_with_reduction_271, multiplication_with_reduction_272, multiplication_with_reduction_273, multiplication_with_reduction_274, multiplication_with_reduction_275, multiplication_with_reduction_276, multiplication_with_reduction_277, multiplication_with_reduction_278, multiplication_with_reduction_279, multiplication_with_reduction_280, multiplication_with_reduction_281, multiplication_with_reduction_282,
-- 0010 multiplication with reduction and prime line equal to 1
multiplication_with_reduction_special_prime_1_0, multiplication_with_reduction_special_prime_1_1,
multiplication_with_reduction_special_prime_1_3, multiplication_with_reduction_special_prime_1_4, multiplication_with_reduction_special_prime_1_5, multiplication_with_reduction_special_prime_1_6, multiplication_with_reduction_special_prime_1_7, multiplication_with_reduction_special_prime_1_8,
multiplication_with_reduction_special_prime_1_10, multiplication_with_reduction_special_prime_1_11, multiplication_with_reduction_special_prime_1_12, multiplication_with_reduction_special_prime_1_13, multiplication_with_reduction_special_prime_1_14, multiplication_with_reduction_special_prime_1_15, multiplication_with_reduction_special_prime_1_16, multiplication_with_reduction_special_prime_1_17, multiplication_with_reduction_special_prime_1_18, multiplication_with_reduction_special_prime_1_19, multiplication_with_reduction_special_prime_1_20,multiplication_with_reduction_special_prime_1_21, multiplication_with_reduction_special_prime_1_22, multiplication_with_reduction_special_prime_1_23,
multiplication_with_reduction_special_prime_1_25, multiplication_with_reduction_special_prime_1_26, multiplication_with_reduction_special_prime_1_27, multiplication_with_reduction_special_prime_1_28, multiplication_with_reduction_special_prime_1_29, multiplication_with_reduction_special_prime_1_30, multiplication_with_reduction_special_prime_1_31, multiplication_with_reduction_special_prime_1_32, multiplication_with_reduction_special_prime_1_33, multiplication_with_reduction_special_prime_1_34, multiplication_with_reduction_special_prime_1_35, multiplication_with_reduction_special_prime_1_36, multiplication_with_reduction_special_prime_1_37, multiplication_with_reduction_special_prime_1_38, multiplication_with_reduction_special_prime_1_39, multiplication_with_reduction_special_prime_1_40, multiplication_with_reduction_special_prime_1_41, multiplication_with_reduction_special_prime_1_42, multiplication_with_reduction_special_prime_1_43, multiplication_with_reduction_special_prime_1_44, multiplication_with_reduction_special_prime_1_45, 
multiplication_with_reduction_special_prime_1_47, multiplication_with_reduction_special_prime_1_48, multiplication_with_reduction_special_prime_1_49, multiplication_with_reduction_special_prime_1_50, multiplication_with_reduction_special_prime_1_51, multiplication_with_reduction_special_prime_1_52, multiplication_with_reduction_special_prime_1_53, multiplication_with_reduction_special_prime_1_54, multiplication_with_reduction_special_prime_1_55, multiplication_with_reduction_special_prime_1_56, multiplication_with_reduction_special_prime_1_57, multiplication_with_reduction_special_prime_1_58, multiplication_with_reduction_special_prime_1_59, multiplication_with_reduction_special_prime_1_60, multiplication_with_reduction_special_prime_1_61, multiplication_with_reduction_special_prime_1_62, multiplication_with_reduction_special_prime_1_63, multiplication_with_reduction_special_prime_1_64, multiplication_with_reduction_special_prime_1_65, multiplication_with_reduction_special_prime_1_66, multiplication_with_reduction_special_prime_1_67, multiplication_with_reduction_special_prime_1_68, multiplication_with_reduction_special_prime_1_69, multiplication_with_reduction_special_prime_1_70, multiplication_with_reduction_special_prime_1_71, multiplication_with_reduction_special_prime_1_72, multiplication_with_reduction_special_prime_1_73, multiplication_with_reduction_special_prime_1_74, multiplication_with_reduction_special_prime_1_75, multiplication_with_reduction_special_prime_1_76, multiplication_with_reduction_special_prime_1_77,
multiplication_with_reduction_special_prime_1_79, multiplication_with_reduction_special_prime_1_80, multiplication_with_reduction_special_prime_1_81, multiplication_with_reduction_special_prime_1_82, multiplication_with_reduction_special_prime_1_83, multiplication_with_reduction_special_prime_1_84, multiplication_with_reduction_special_prime_1_85, multiplication_with_reduction_special_prime_1_86, multiplication_with_reduction_special_prime_1_87, multiplication_with_reduction_special_prime_1_88, multiplication_with_reduction_special_prime_1_89, multiplication_with_reduction_special_prime_1_90,
multiplication_with_reduction_special_prime_1_91, multiplication_with_reduction_special_prime_1_92, multiplication_with_reduction_special_prime_1_93, multiplication_with_reduction_special_prime_1_94, multiplication_with_reduction_special_prime_1_95, multiplication_with_reduction_special_prime_1_96, multiplication_with_reduction_special_prime_1_97, multiplication_with_reduction_special_prime_1_98, multiplication_with_reduction_special_prime_1_99, multiplication_with_reduction_special_prime_1_100, multiplication_with_reduction_special_prime_1_101, multiplication_with_reduction_special_prime_1_102, multiplication_with_reduction_special_prime_1_103, multiplication_with_reduction_special_prime_1_104, multiplication_with_reduction_special_prime_1_105, multiplication_with_reduction_special_prime_1_106, multiplication_with_reduction_special_prime_1_107, multiplication_with_reduction_special_prime_1_108, multiplication_with_reduction_special_prime_1_109, multiplication_with_reduction_special_prime_1_110, multiplication_with_reduction_special_prime_1_111, multiplication_with_reduction_special_prime_1_112, multiplication_with_reduction_special_prime_1_113, multiplication_with_reduction_special_prime_1_114, multiplication_with_reduction_special_prime_1_115, multiplication_with_reduction_special_prime_1_116, multiplication_with_reduction_special_prime_1_117, multiplication_with_reduction_special_prime_1_118, multiplication_with_reduction_special_prime_1_119, multiplication_with_reduction_special_prime_1_120, multiplication_with_reduction_special_prime_1_121, 
multiplication_with_reduction_special_prime_1_123, multiplication_with_reduction_special_prime_1_124, multiplication_with_reduction_special_prime_1_125, multiplication_with_reduction_special_prime_1_126, multiplication_with_reduction_special_prime_1_127, multiplication_with_reduction_special_prime_1_128, multiplication_with_reduction_special_prime_1_129, multiplication_with_reduction_special_prime_1_130, multiplication_with_reduction_special_prime_1_131, multiplication_with_reduction_special_prime_1_132, multiplication_with_reduction_special_prime_1_133, multiplication_with_reduction_special_prime_1_134, multiplication_with_reduction_special_prime_1_135, multiplication_with_reduction_special_prime_1_136, multiplication_with_reduction_special_prime_1_137, multiplication_with_reduction_special_prime_1_138, multiplication_with_reduction_special_prime_1_139, multiplication_with_reduction_special_prime_1_140, multiplication_with_reduction_special_prime_1_141, multiplication_with_reduction_special_prime_1_142, multiplication_with_reduction_special_prime_1_143, multiplication_with_reduction_special_prime_1_144, multiplication_with_reduction_special_prime_1_145, multiplication_with_reduction_special_prime_1_146, multiplication_with_reduction_special_prime_1_147, multiplication_with_reduction_special_prime_1_148, multiplication_with_reduction_special_prime_1_149, multiplication_with_reduction_special_prime_1_150, multiplication_with_reduction_special_prime_1_151, multiplication_with_reduction_special_prime_1_152, multiplication_with_reduction_special_prime_1_153, multiplication_with_reduction_special_prime_1_154, multiplication_with_reduction_special_prime_1_155, multiplication_with_reduction_special_prime_1_156, multiplication_with_reduction_special_prime_1_157, multiplication_with_reduction_special_prime_1_158, multiplication_with_reduction_special_prime_1_159, multiplication_with_reduction_special_prime_1_160, multiplication_with_reduction_special_prime_1_161, multiplication_with_reduction_special_prime_1_162, multiplication_with_reduction_special_prime_1_163, multiplication_with_reduction_special_prime_1_164, multiplication_with_reduction_special_prime_1_165, multiplication_with_reduction_special_prime_1_166, multiplication_with_reduction_special_prime_1_167, multiplication_with_reduction_special_prime_1_168, multiplication_with_reduction_special_prime_1_169, multiplication_with_reduction_special_prime_1_170, multiplication_with_reduction_special_prime_1_171, multiplication_with_reduction_special_prime_1_172, multiplication_with_reduction_special_prime_1_173, multiplication_with_reduction_special_prime_1_174, multiplication_with_reduction_special_prime_1_175, multiplication_with_reduction_special_prime_1_176, multiplication_with_reduction_special_prime_1_177, multiplication_with_reduction_special_prime_1_178, multiplication_with_reduction_special_prime_1_179,
multiplication_with_reduction_special_prime_1_181, multiplication_with_reduction_special_prime_1_182, multiplication_with_reduction_special_prime_1_183, multiplication_with_reduction_special_prime_1_184, multiplication_with_reduction_special_prime_1_185, multiplication_with_reduction_special_prime_1_186, multiplication_with_reduction_special_prime_1_187, multiplication_with_reduction_special_prime_1_188, multiplication_with_reduction_special_prime_1_189, multiplication_with_reduction_special_prime_1_190, multiplication_with_reduction_special_prime_1_191, multiplication_with_reduction_special_prime_1_192, multiplication_with_reduction_special_prime_1_193, multiplication_with_reduction_special_prime_1_194, multiplication_with_reduction_special_prime_1_195, multiplication_with_reduction_special_prime_1_196, multiplication_with_reduction_special_prime_1_197, multiplication_with_reduction_special_prime_1_198, multiplication_with_reduction_special_prime_1_199, multiplication_with_reduction_special_prime_1_200, multiplication_with_reduction_special_prime_1_201, multiplication_with_reduction_special_prime_1_202, multiplication_with_reduction_special_prime_1_203, multiplication_with_reduction_special_prime_1_204, multiplication_with_reduction_special_prime_1_205, multiplication_with_reduction_special_prime_1_206, multiplication_with_reduction_special_prime_1_207, multiplication_with_reduction_special_prime_1_208, multiplication_with_reduction_special_prime_1_209, multiplication_with_reduction_special_prime_1_210, multiplication_with_reduction_special_prime_1_211, multiplication_with_reduction_special_prime_1_212, multiplication_with_reduction_special_prime_1_213, multiplication_with_reduction_special_prime_1_214, multiplication_with_reduction_special_prime_1_215, multiplication_with_reduction_special_prime_1_216, multiplication_with_reduction_special_prime_1_217, multiplication_with_reduction_special_prime_1_218, multiplication_with_reduction_special_prime_1_219, multiplication_with_reduction_special_prime_1_220, multiplication_with_reduction_special_prime_1_221, multiplication_with_reduction_special_prime_1_222, multiplication_with_reduction_special_prime_1_223, multiplication_with_reduction_special_prime_1_224, multiplication_with_reduction_special_prime_1_225, multiplication_with_reduction_special_prime_1_226, multiplication_with_reduction_special_prime_1_227, multiplication_with_reduction_special_prime_1_228, multiplication_with_reduction_special_prime_1_229, multiplication_with_reduction_special_prime_1_230, multiplication_with_reduction_special_prime_1_231, multiplication_with_reduction_special_prime_1_232, multiplication_with_reduction_special_prime_1_233, multiplication_with_reduction_special_prime_1_234, multiplication_with_reduction_special_prime_1_235, multiplication_with_reduction_special_prime_1_236, multiplication_with_reduction_special_prime_1_237, multiplication_with_reduction_special_prime_1_238, multiplication_with_reduction_special_prime_1_239, multiplication_with_reduction_special_prime_1_240, multiplication_with_reduction_special_prime_1_241, multiplication_with_reduction_special_prime_1_242, multiplication_with_reduction_special_prime_1_243, multiplication_with_reduction_special_prime_1_244, multiplication_with_reduction_special_prime_1_245, multiplication_with_reduction_special_prime_1_246, multiplication_with_reduction_special_prime_1_247, multiplication_with_reduction_special_prime_1_248, multiplication_with_reduction_special_prime_1_249, multiplication_with_reduction_special_prime_1_250, multiplication_with_reduction_special_prime_1_251, multiplication_with_reduction_special_prime_1_252, multiplication_with_reduction_special_prime_1_253,
multiplication_with_reduction_special_prime_2_0, multiplication_with_reduction_special_prime_2_1, multiplication_with_reduction_special_prime_2_2, multiplication_with_reduction_special_prime_2_3,
multiplication_with_reduction_special_prime_2_5, multiplication_with_reduction_special_prime_2_6, multiplication_with_reduction_special_prime_2_7, multiplication_with_reduction_special_prime_2_8, multiplication_with_reduction_special_prime_2_9, multiplication_with_reduction_special_prime_2_10, multiplication_with_reduction_special_prime_2_11, multiplication_with_reduction_special_prime_2_12, multiplication_with_reduction_special_prime_2_13, multiplication_with_reduction_special_prime_2_14, multiplication_with_reduction_special_prime_2_15,
multiplication_with_reduction_special_prime_2_17, multiplication_with_reduction_special_prime_2_18, multiplication_with_reduction_special_prime_2_19, multiplication_with_reduction_special_prime_2_20, multiplication_with_reduction_special_prime_2_21, multiplication_with_reduction_special_prime_2_22, multiplication_with_reduction_special_prime_2_23, multiplication_with_reduction_special_prime_2_24, multiplication_with_reduction_special_prime_2_25, multiplication_with_reduction_special_prime_2_26, multiplication_with_reduction_special_prime_2_27, multiplication_with_reduction_special_prime_2_28, multiplication_with_reduction_special_prime_2_29, multiplication_with_reduction_special_prime_2_30, multiplication_with_reduction_special_prime_2_31, multiplication_with_reduction_special_prime_2_32, multiplication_with_reduction_special_prime_2_33, multiplication_with_reduction_special_prime_2_34, multiplication_with_reduction_special_prime_2_35,
multiplication_with_reduction_special_prime_2_37, multiplication_with_reduction_special_prime_2_38, multiplication_with_reduction_special_prime_2_39, multiplication_with_reduction_special_prime_2_40, multiplication_with_reduction_special_prime_2_41, multiplication_with_reduction_special_prime_2_42, multiplication_with_reduction_special_prime_2_43, multiplication_with_reduction_special_prime_2_44, multiplication_with_reduction_special_prime_2_45, multiplication_with_reduction_special_prime_2_46, multiplication_with_reduction_special_prime_2_47, multiplication_with_reduction_special_prime_2_48, multiplication_with_reduction_special_prime_2_49, multiplication_with_reduction_special_prime_2_50, multiplication_with_reduction_special_prime_2_51, multiplication_with_reduction_special_prime_2_52, multiplication_with_reduction_special_prime_2_53, multiplication_with_reduction_special_prime_2_54, multiplication_with_reduction_special_prime_2_55, multiplication_with_reduction_special_prime_2_56, multiplication_with_reduction_special_prime_2_57, multiplication_with_reduction_special_prime_2_58, multiplication_with_reduction_special_prime_2_59, multiplication_with_reduction_special_prime_2_60, multiplication_with_reduction_special_prime_2_61, multiplication_with_reduction_special_prime_2_62, multiplication_with_reduction_special_prime_2_63, multiplication_with_reduction_special_prime_2_64, multiplication_with_reduction_special_prime_2_65,
multiplication_with_reduction_special_prime_2_67, multiplication_with_reduction_special_prime_2_68, multiplication_with_reduction_special_prime_2_69, multiplication_with_reduction_special_prime_2_70, multiplication_with_reduction_special_prime_2_71, multiplication_with_reduction_special_prime_2_72, multiplication_with_reduction_special_prime_2_73, multiplication_with_reduction_special_prime_2_74, multiplication_with_reduction_special_prime_2_75, multiplication_with_reduction_special_prime_2_76, multiplication_with_reduction_special_prime_2_77, multiplication_with_reduction_special_prime_2_78, multiplication_with_reduction_special_prime_2_79, multiplication_with_reduction_special_prime_2_80, multiplication_with_reduction_special_prime_2_81, multiplication_with_reduction_special_prime_2_82, multiplication_with_reduction_special_prime_2_83, multiplication_with_reduction_special_prime_2_84, multiplication_with_reduction_special_prime_2_85, multiplication_with_reduction_special_prime_2_86, multiplication_with_reduction_special_prime_2_87, multiplication_with_reduction_special_prime_2_88, multiplication_with_reduction_special_prime_2_89, multiplication_with_reduction_special_prime_2_90, multiplication_with_reduction_special_prime_2_91, multiplication_with_reduction_special_prime_2_92, multiplication_with_reduction_special_prime_2_93, multiplication_with_reduction_special_prime_2_94, multiplication_with_reduction_special_prime_2_95, multiplication_with_reduction_special_prime_2_96, multiplication_with_reduction_special_prime_2_97, multiplication_with_reduction_special_prime_2_98, multiplication_with_reduction_special_prime_2_99, multiplication_with_reduction_special_prime_2_100, multiplication_with_reduction_special_prime_2_101, multiplication_with_reduction_special_prime_2_102, multiplication_with_reduction_special_prime_2_103, multiplication_with_reduction_special_prime_2_104, multiplication_with_reduction_special_prime_2_105, multiplication_with_reduction_special_prime_2_106, multiplication_with_reduction_special_prime_2_107,
multiplication_with_reduction_special_prime_2_109, multiplication_with_reduction_special_prime_2_110, multiplication_with_reduction_special_prime_2_111, multiplication_with_reduction_special_prime_2_112, multiplication_with_reduction_special_prime_2_113, multiplication_with_reduction_special_prime_2_114, multiplication_with_reduction_special_prime_2_115, multiplication_with_reduction_special_prime_2_116, multiplication_with_reduction_special_prime_2_117, multiplication_with_reduction_special_prime_2_118, multiplication_with_reduction_special_prime_2_119, multiplication_with_reduction_special_prime_2_120, multiplication_with_reduction_special_prime_2_121, multiplication_with_reduction_special_prime_2_122, multiplication_with_reduction_special_prime_2_123, multiplication_with_reduction_special_prime_2_124, multiplication_with_reduction_special_prime_2_125, multiplication_with_reduction_special_prime_2_126, multiplication_with_reduction_special_prime_2_127, multiplication_with_reduction_special_prime_2_128, multiplication_with_reduction_special_prime_2_129, multiplication_with_reduction_special_prime_2_130, multiplication_with_reduction_special_prime_2_131, multiplication_with_reduction_special_prime_2_132, multiplication_with_reduction_special_prime_2_133, multiplication_with_reduction_special_prime_2_134, multiplication_with_reduction_special_prime_2_135, multiplication_with_reduction_special_prime_2_136, multiplication_with_reduction_special_prime_2_137, multiplication_with_reduction_special_prime_2_138, multiplication_with_reduction_special_prime_2_139, multiplication_with_reduction_special_prime_2_140, multiplication_with_reduction_special_prime_2_141, multiplication_with_reduction_special_prime_2_142, multiplication_with_reduction_special_prime_2_143, multiplication_with_reduction_special_prime_2_144, multiplication_with_reduction_special_prime_2_145, multiplication_with_reduction_special_prime_2_146, multiplication_with_reduction_special_prime_2_147, multiplication_with_reduction_special_prime_2_148, multiplication_with_reduction_special_prime_2_149, multiplication_with_reduction_special_prime_2_150, multiplication_with_reduction_special_prime_2_151, multiplication_with_reduction_special_prime_2_152, multiplication_with_reduction_special_prime_2_153, multiplication_with_reduction_special_prime_2_154, multiplication_with_reduction_special_prime_2_155, multiplication_with_reduction_special_prime_2_156, multiplication_with_reduction_special_prime_2_157, multiplication_with_reduction_special_prime_2_158, multiplication_with_reduction_special_prime_2_159, multiplication_with_reduction_special_prime_2_160, multiplication_with_reduction_special_prime_2_161, multiplication_with_reduction_special_prime_2_162, multiplication_with_reduction_special_prime_2_163,
multiplication_with_reduction_special_prime_2_165, multiplication_with_reduction_special_prime_2_166, multiplication_with_reduction_special_prime_2_167, multiplication_with_reduction_special_prime_2_168, multiplication_with_reduction_special_prime_2_169, multiplication_with_reduction_special_prime_2_170, multiplication_with_reduction_special_prime_2_171, multiplication_with_reduction_special_prime_2_172, multiplication_with_reduction_special_prime_2_173, multiplication_with_reduction_special_prime_2_174, multiplication_with_reduction_special_prime_2_175, multiplication_with_reduction_special_prime_2_176, multiplication_with_reduction_special_prime_2_177, multiplication_with_reduction_special_prime_2_178, multiplication_with_reduction_special_prime_2_179, multiplication_with_reduction_special_prime_2_180, multiplication_with_reduction_special_prime_2_181, multiplication_with_reduction_special_prime_2_182, multiplication_with_reduction_special_prime_2_183, multiplication_with_reduction_special_prime_2_184, multiplication_with_reduction_special_prime_2_185, multiplication_with_reduction_special_prime_2_186, multiplication_with_reduction_special_prime_2_187, multiplication_with_reduction_special_prime_2_188, multiplication_with_reduction_special_prime_2_189, multiplication_with_reduction_special_prime_2_190, multiplication_with_reduction_special_prime_2_191, multiplication_with_reduction_special_prime_2_192, multiplication_with_reduction_special_prime_2_193, multiplication_with_reduction_special_prime_2_194, multiplication_with_reduction_special_prime_2_195, multiplication_with_reduction_special_prime_2_196, multiplication_with_reduction_special_prime_2_197, multiplication_with_reduction_special_prime_2_198, multiplication_with_reduction_special_prime_2_199, multiplication_with_reduction_special_prime_2_200, multiplication_with_reduction_special_prime_2_201, multiplication_with_reduction_special_prime_2_202, multiplication_with_reduction_special_prime_2_203, multiplication_with_reduction_special_prime_2_204, multiplication_with_reduction_special_prime_2_205, multiplication_with_reduction_special_prime_2_206, multiplication_with_reduction_special_prime_2_207, multiplication_with_reduction_special_prime_2_208, multiplication_with_reduction_special_prime_2_209, multiplication_with_reduction_special_prime_2_210, multiplication_with_reduction_special_prime_2_211, multiplication_with_reduction_special_prime_2_212, multiplication_with_reduction_special_prime_2_213, multiplication_with_reduction_special_prime_2_214, multiplication_with_reduction_special_prime_2_215, multiplication_with_reduction_special_prime_2_216, multiplication_with_reduction_special_prime_2_217, multiplication_with_reduction_special_prime_2_218, multiplication_with_reduction_special_prime_2_219, multiplication_with_reduction_special_prime_2_220, multiplication_with_reduction_special_prime_2_221, multiplication_with_reduction_special_prime_2_222, multiplication_with_reduction_special_prime_2_223, multiplication_with_reduction_special_prime_2_224, multiplication_with_reduction_special_prime_2_225, multiplication_with_reduction_special_prime_2_226, multiplication_with_reduction_special_prime_2_227, multiplication_with_reduction_special_prime_2_228, multiplication_with_reduction_special_prime_2_229, multiplication_with_reduction_special_prime_2_230, multiplication_with_reduction_special_prime_2_231, multiplication_with_reduction_special_prime_2_232, multiplication_with_reduction_special_prime_2_233, multiplication_with_reduction_special_prime_2_234, multiplication_with_reduction_special_prime_2_235,
multiplication_with_reduction_special_prime_3_0, multiplication_with_reduction_special_prime_3_1, multiplication_with_reduction_special_prime_3_2, multiplication_with_reduction_special_prime_3_3, multiplication_with_reduction_special_prime_3_4, multiplication_with_reduction_special_prime_3_5, multiplication_with_reduction_special_prime_3_6, multiplication_with_reduction_special_prime_3_7, multiplication_with_reduction_special_prime_3_8, 
multiplication_with_reduction_special_prime_3_10, multiplication_with_reduction_special_prime_3_11, multiplication_with_reduction_special_prime_3_12, multiplication_with_reduction_special_prime_3_13, multiplication_with_reduction_special_prime_3_14, multiplication_with_reduction_special_prime_3_15, multiplication_with_reduction_special_prime_3_16, multiplication_with_reduction_special_prime_3_17, multiplication_with_reduction_special_prime_3_18, multiplication_with_reduction_special_prime_3_19, multiplication_with_reduction_special_prime_3_20, multiplication_with_reduction_special_prime_3_21, multiplication_with_reduction_special_prime_3_22, multiplication_with_reduction_special_prime_3_23, multiplication_with_reduction_special_prime_3_24, multiplication_with_reduction_special_prime_3_25,
multiplication_with_reduction_special_prime_3_27, multiplication_with_reduction_special_prime_3_28, multiplication_with_reduction_special_prime_3_29, multiplication_with_reduction_special_prime_3_30, multiplication_with_reduction_special_prime_3_31, multiplication_with_reduction_special_prime_3_32, multiplication_with_reduction_special_prime_3_33, multiplication_with_reduction_special_prime_3_34, multiplication_with_reduction_special_prime_3_35, multiplication_with_reduction_special_prime_3_36, multiplication_with_reduction_special_prime_3_37, multiplication_with_reduction_special_prime_3_38, multiplication_with_reduction_special_prime_3_39, multiplication_with_reduction_special_prime_3_40, multiplication_with_reduction_special_prime_3_41, multiplication_with_reduction_special_prime_3_42, multiplication_with_reduction_special_prime_3_43, multiplication_with_reduction_special_prime_3_44, multiplication_with_reduction_special_prime_3_45, multiplication_with_reduction_special_prime_3_46, multiplication_with_reduction_special_prime_3_47, multiplication_with_reduction_special_prime_3_48, multiplication_with_reduction_special_prime_3_49, multiplication_with_reduction_special_prime_3_50, multiplication_with_reduction_special_prime_3_51, multiplication_with_reduction_special_prime_3_52,
multiplication_with_reduction_special_prime_3_54, multiplication_with_reduction_special_prime_3_55, multiplication_with_reduction_special_prime_3_56, multiplication_with_reduction_special_prime_3_57, multiplication_with_reduction_special_prime_3_58, multiplication_with_reduction_special_prime_3_59, multiplication_with_reduction_special_prime_3_60, multiplication_with_reduction_special_prime_3_61, multiplication_with_reduction_special_prime_3_62, multiplication_with_reduction_special_prime_3_63, multiplication_with_reduction_special_prime_3_64, multiplication_with_reduction_special_prime_3_65, multiplication_with_reduction_special_prime_3_66, multiplication_with_reduction_special_prime_3_67, multiplication_with_reduction_special_prime_3_68, multiplication_with_reduction_special_prime_3_69, multiplication_with_reduction_special_prime_3_70, multiplication_with_reduction_special_prime_3_71, multiplication_with_reduction_special_prime_3_72, multiplication_with_reduction_special_prime_3_73, multiplication_with_reduction_special_prime_3_74, multiplication_with_reduction_special_prime_3_75, multiplication_with_reduction_special_prime_3_76, multiplication_with_reduction_special_prime_3_77, multiplication_with_reduction_special_prime_3_78, multiplication_with_reduction_special_prime_3_79, multiplication_with_reduction_special_prime_3_80, multiplication_with_reduction_special_prime_3_81, multiplication_with_reduction_special_prime_3_82, multiplication_with_reduction_special_prime_3_83, multiplication_with_reduction_special_prime_3_84, multiplication_with_reduction_special_prime_3_85, multiplication_with_reduction_special_prime_3_86, multiplication_with_reduction_special_prime_3_87, multiplication_with_reduction_special_prime_3_88, multiplication_with_reduction_special_prime_3_89, multiplication_with_reduction_special_prime_3_90, multiplication_with_reduction_special_prime_3_91,
multiplication_with_reduction_special_prime_3_93, multiplication_with_reduction_special_prime_3_94, multiplication_with_reduction_special_prime_3_95, multiplication_with_reduction_special_prime_3_96, multiplication_with_reduction_special_prime_3_97, multiplication_with_reduction_special_prime_3_98, multiplication_with_reduction_special_prime_3_99, multiplication_with_reduction_special_prime_3_100, multiplication_with_reduction_special_prime_3_101, multiplication_with_reduction_special_prime_3_102, multiplication_with_reduction_special_prime_3_103, multiplication_with_reduction_special_prime_3_104, multiplication_with_reduction_special_prime_3_105, multiplication_with_reduction_special_prime_3_106, multiplication_with_reduction_special_prime_3_107, multiplication_with_reduction_special_prime_3_108, multiplication_with_reduction_special_prime_3_109, multiplication_with_reduction_special_prime_3_110, multiplication_with_reduction_special_prime_3_111, multiplication_with_reduction_special_prime_3_112, multiplication_with_reduction_special_prime_3_113, multiplication_with_reduction_special_prime_3_114, multiplication_with_reduction_special_prime_3_115, multiplication_with_reduction_special_prime_3_116, multiplication_with_reduction_special_prime_3_117, multiplication_with_reduction_special_prime_3_118, multiplication_with_reduction_special_prime_3_119, multiplication_with_reduction_special_prime_3_120, multiplication_with_reduction_special_prime_3_121, multiplication_with_reduction_special_prime_3_122, multiplication_with_reduction_special_prime_3_123, multiplication_with_reduction_special_prime_3_124, multiplication_with_reduction_special_prime_3_125, multiplication_with_reduction_special_prime_3_126, multiplication_with_reduction_special_prime_3_127, multiplication_with_reduction_special_prime_3_128, multiplication_with_reduction_special_prime_3_129, multiplication_with_reduction_special_prime_3_130, multiplication_with_reduction_special_prime_3_131, multiplication_with_reduction_special_prime_3_132, multiplication_with_reduction_special_prime_3_133, multiplication_with_reduction_special_prime_3_134, multiplication_with_reduction_special_prime_3_135, multiplication_with_reduction_special_prime_3_136, multiplication_with_reduction_special_prime_3_137, multiplication_with_reduction_special_prime_3_138, multiplication_with_reduction_special_prime_3_139, multiplication_with_reduction_special_prime_3_140, multiplication_with_reduction_special_prime_3_141, multiplication_with_reduction_special_prime_3_142, multiplication_with_reduction_special_prime_3_143, multiplication_with_reduction_special_prime_3_144,
multiplication_with_reduction_special_prime_3_146, multiplication_with_reduction_special_prime_3_147, multiplication_with_reduction_special_prime_3_148, multiplication_with_reduction_special_prime_3_149, multiplication_with_reduction_special_prime_3_150, multiplication_with_reduction_special_prime_3_151, multiplication_with_reduction_special_prime_3_152, multiplication_with_reduction_special_prime_3_153, multiplication_with_reduction_special_prime_3_154, multiplication_with_reduction_special_prime_3_155, multiplication_with_reduction_special_prime_3_156, multiplication_with_reduction_special_prime_3_157, multiplication_with_reduction_special_prime_3_158, multiplication_with_reduction_special_prime_3_159, multiplication_with_reduction_special_prime_3_160, multiplication_with_reduction_special_prime_3_161, multiplication_with_reduction_special_prime_3_162, multiplication_with_reduction_special_prime_3_163, multiplication_with_reduction_special_prime_3_164, multiplication_with_reduction_special_prime_3_165, multiplication_with_reduction_special_prime_3_166, multiplication_with_reduction_special_prime_3_167, multiplication_with_reduction_special_prime_3_168, multiplication_with_reduction_special_prime_3_169, multiplication_with_reduction_special_prime_3_170, multiplication_with_reduction_special_prime_3_171, multiplication_with_reduction_special_prime_3_172, multiplication_with_reduction_special_prime_3_173, multiplication_with_reduction_special_prime_3_174, multiplication_with_reduction_special_prime_3_175, multiplication_with_reduction_special_prime_3_176, multiplication_with_reduction_special_prime_3_177, multiplication_with_reduction_special_prime_3_178, multiplication_with_reduction_special_prime_3_179, multiplication_with_reduction_special_prime_3_180, multiplication_with_reduction_special_prime_3_181, multiplication_with_reduction_special_prime_3_182, multiplication_with_reduction_special_prime_3_183, multiplication_with_reduction_special_prime_3_184, multiplication_with_reduction_special_prime_3_185, multiplication_with_reduction_special_prime_3_186, multiplication_with_reduction_special_prime_3_187, multiplication_with_reduction_special_prime_3_188, multiplication_with_reduction_special_prime_3_189, multiplication_with_reduction_special_prime_3_190, multiplication_with_reduction_special_prime_3_191, multiplication_with_reduction_special_prime_3_192, multiplication_with_reduction_special_prime_3_193, multiplication_with_reduction_special_prime_3_194, multiplication_with_reduction_special_prime_3_195, multiplication_with_reduction_special_prime_3_196, multiplication_with_reduction_special_prime_3_197, multiplication_with_reduction_special_prime_3_198, multiplication_with_reduction_special_prime_3_199, multiplication_with_reduction_special_prime_3_200, multiplication_with_reduction_special_prime_3_201, multiplication_with_reduction_special_prime_3_202, multiplication_with_reduction_special_prime_3_203, multiplication_with_reduction_special_prime_3_204, multiplication_with_reduction_special_prime_3_205, multiplication_with_reduction_special_prime_3_206, multiplication_with_reduction_special_prime_3_207, multiplication_with_reduction_special_prime_3_208, multiplication_with_reduction_special_prime_3_209, multiplication_with_reduction_special_prime_3_210, multiplication_with_reduction_special_prime_3_211, multiplication_with_reduction_special_prime_3_212, multiplication_with_reduction_special_prime_3_213,
-- 0011 square with reduction and prime line not equal to 1
square_with_reduction_0, square_with_reduction_1, square_with_reduction_2, square_with_reduction_3,
square_with_reduction_5, square_with_reduction_6, square_with_reduction_7, square_with_reduction_8, square_with_reduction_9, square_with_reduction_10, square_with_reduction_11, square_with_reduction_12, square_with_reduction_13,
square_with_reduction_15, square_with_reduction_16, square_with_reduction_17, square_with_reduction_18, square_with_reduction_19, square_with_reduction_20, square_with_reduction_21, square_with_reduction_22, square_with_reduction_23, square_with_reduction_24, square_with_reduction_25, square_with_reduction_26, square_with_reduction_27, square_with_reduction_28, 
square_with_reduction_30, square_with_reduction_31, square_with_reduction_32, square_with_reduction_33, square_with_reduction_34, square_with_reduction_35, square_with_reduction_36, square_with_reduction_37, square_with_reduction_38, square_with_reduction_39, square_with_reduction_40, square_with_reduction_41, square_with_reduction_42, square_with_reduction_43, square_with_reduction_44, square_with_reduction_45, square_with_reduction_46, square_with_reduction_47, square_with_reduction_48, square_with_reduction_49,
square_with_reduction_51, square_with_reduction_52, square_with_reduction_53, square_with_reduction_54, square_with_reduction_55, square_with_reduction_56, square_with_reduction_57, square_with_reduction_58, square_with_reduction_59, square_with_reduction_60, square_with_reduction_61, square_with_reduction_62, square_with_reduction_63, square_with_reduction_64, square_with_reduction_65, square_with_reduction_66, square_with_reduction_67, square_with_reduction_68, square_with_reduction_69, square_with_reduction_70, square_with_reduction_71, square_with_reduction_72, square_with_reduction_73, square_with_reduction_74, square_with_reduction_75, square_with_reduction_76, square_with_reduction_77, square_with_reduction_78,
square_with_reduction_80, square_with_reduction_81, square_with_reduction_82, square_with_reduction_83, square_with_reduction_84, square_with_reduction_85, square_with_reduction_86, square_with_reduction_87, square_with_reduction_88, square_with_reduction_89, square_with_reduction_90, square_with_reduction_91, square_with_reduction_92, square_with_reduction_93, square_with_reduction_94, square_with_reduction_95, square_with_reduction_96, square_with_reduction_97, square_with_reduction_98, square_with_reduction_99, square_with_reduction_100, square_with_reduction_101, square_with_reduction_102, square_with_reduction_103, square_with_reduction_104, square_with_reduction_105, square_with_reduction_106, square_with_reduction_107, square_with_reduction_108, square_with_reduction_109, square_with_reduction_110, square_with_reduction_111, square_with_reduction_112, square_with_reduction_113, square_with_reduction_114, square_with_reduction_115, square_with_reduction_116,
square_with_reduction_118, square_with_reduction_119, square_with_reduction_120, square_with_reduction_121, square_with_reduction_122, square_with_reduction_123, square_with_reduction_124, square_with_reduction_125, square_with_reduction_126, square_with_reduction_127, square_with_reduction_128, square_with_reduction_129, square_with_reduction_130, square_with_reduction_131, square_with_reduction_132, square_with_reduction_133, square_with_reduction_134, square_with_reduction_135, square_with_reduction_136, square_with_reduction_137, square_with_reduction_138, square_with_reduction_139, square_with_reduction_140, square_with_reduction_141, square_with_reduction_142, square_with_reduction_143, square_with_reduction_144, square_with_reduction_145, square_with_reduction_146, square_with_reduction_147, square_with_reduction_148, square_with_reduction_149, square_with_reduction_150, square_with_reduction_151, square_with_reduction_152, square_with_reduction_153, square_with_reduction_154, square_with_reduction_155, square_with_reduction_156, square_with_reduction_157, square_with_reduction_158, square_with_reduction_159, square_with_reduction_160, square_with_reduction_161, square_with_reduction_162, square_with_reduction_163, square_with_reduction_164, square_with_reduction_165,
square_with_reduction_167, square_with_reduction_168, square_with_reduction_169, square_with_reduction_170, square_with_reduction_171, square_with_reduction_172, square_with_reduction_173, square_with_reduction_174, square_with_reduction_175, square_with_reduction_176, square_with_reduction_177, square_with_reduction_178, square_with_reduction_179, square_with_reduction_180, square_with_reduction_181, square_with_reduction_182, square_with_reduction_183, square_with_reduction_184, square_with_reduction_185, square_with_reduction_186, square_with_reduction_187, square_with_reduction_188, square_with_reduction_189, square_with_reduction_190, square_with_reduction_191, square_with_reduction_192, square_with_reduction_193, square_with_reduction_194, square_with_reduction_195, square_with_reduction_196, square_with_reduction_197, square_with_reduction_198, square_with_reduction_199, square_with_reduction_200, square_with_reduction_201, square_with_reduction_202, square_with_reduction_203, square_with_reduction_204, square_with_reduction_205, square_with_reduction_206, square_with_reduction_207, square_with_reduction_208, square_with_reduction_209, square_with_reduction_210, square_with_reduction_211, square_with_reduction_212, square_with_reduction_213, square_with_reduction_214, square_with_reduction_215, square_with_reduction_216, square_with_reduction_217, square_with_reduction_218, square_with_reduction_219, square_with_reduction_220, square_with_reduction_221, square_with_reduction_222, square_with_reduction_223, square_with_reduction_224, square_with_reduction_225, square_with_reduction_226,
-- 0011 square with reduction and prime line equal to 1
square_with_reduction_special_prime_1_0, square_with_reduction_special_prime_1_1,
square_with_reduction_special_prime_1_3, square_with_reduction_special_prime_1_4, square_with_reduction_special_prime_1_5, square_with_reduction_special_prime_1_6, square_with_reduction_special_prime_1_7,
square_with_reduction_special_prime_1_9, square_with_reduction_special_prime_1_10, square_with_reduction_special_prime_1_11, square_with_reduction_special_prime_1_12, square_with_reduction_special_prime_1_13, square_with_reduction_special_prime_1_14, square_with_reduction_special_prime_1_15, square_with_reduction_special_prime_1_16, square_with_reduction_special_prime_1_17, square_with_reduction_special_prime_1_18,
square_with_reduction_special_prime_1_20, square_with_reduction_special_prime_1_21, square_with_reduction_special_prime_1_22, square_with_reduction_special_prime_1_23, square_with_reduction_special_prime_1_24, square_with_reduction_special_prime_1_25, square_with_reduction_special_prime_1_26, square_with_reduction_special_prime_1_27, square_with_reduction_special_prime_1_28, square_with_reduction_special_prime_1_29, square_with_reduction_special_prime_1_30, square_with_reduction_special_prime_1_31, square_with_reduction_special_prime_1_32, square_with_reduction_special_prime_1_33, square_with_reduction_special_prime_1_34, square_with_reduction_special_prime_1_35,
square_with_reduction_special_prime_1_37, square_with_reduction_special_prime_1_38, square_with_reduction_special_prime_1_39, square_with_reduction_special_prime_1_40, square_with_reduction_special_prime_1_41, square_with_reduction_special_prime_1_42, square_with_reduction_special_prime_1_43, square_with_reduction_special_prime_1_44, square_with_reduction_special_prime_1_45, square_with_reduction_special_prime_1_46, square_with_reduction_special_prime_1_47, square_with_reduction_special_prime_1_48, square_with_reduction_special_prime_1_49, square_with_reduction_special_prime_1_50, square_with_reduction_special_prime_1_51, square_with_reduction_special_prime_1_52, square_with_reduction_special_prime_1_53, square_with_reduction_special_prime_1_54, square_with_reduction_special_prime_1_55, square_with_reduction_special_prime_1_56, square_with_reduction_special_prime_1_57, square_with_reduction_special_prime_1_58, square_with_reduction_special_prime_1_59, square_with_reduction_special_prime_1_60, 
square_with_reduction_special_prime_1_62, square_with_reduction_special_prime_1_63, square_with_reduction_special_prime_1_64, square_with_reduction_special_prime_1_65, square_with_reduction_special_prime_1_66, square_with_reduction_special_prime_1_67, square_with_reduction_special_prime_1_68, square_with_reduction_special_prime_1_69, square_with_reduction_special_prime_1_70, square_with_reduction_special_prime_1_71, square_with_reduction_special_prime_1_72, square_with_reduction_special_prime_1_73, square_with_reduction_special_prime_1_74, square_with_reduction_special_prime_1_75, square_with_reduction_special_prime_1_76, square_with_reduction_special_prime_1_77, square_with_reduction_special_prime_1_78, square_with_reduction_special_prime_1_79, square_with_reduction_special_prime_1_80, square_with_reduction_special_prime_1_81, square_with_reduction_special_prime_1_82, square_with_reduction_special_prime_1_83, square_with_reduction_special_prime_1_84, square_with_reduction_special_prime_1_85, square_with_reduction_special_prime_1_86, square_with_reduction_special_prime_1_87, square_with_reduction_special_prime_1_88, square_with_reduction_special_prime_1_89, square_with_reduction_special_prime_1_90, square_with_reduction_special_prime_1_91, square_with_reduction_special_prime_1_92, square_with_reduction_special_prime_1_93, square_with_reduction_special_prime_1_94, 
square_with_reduction_special_prime_1_96, square_with_reduction_special_prime_1_97, square_with_reduction_special_prime_1_98, square_with_reduction_special_prime_1_99, square_with_reduction_special_prime_1_100, square_with_reduction_special_prime_1_101, square_with_reduction_special_prime_1_102, square_with_reduction_special_prime_1_103, square_with_reduction_special_prime_1_104, square_with_reduction_special_prime_1_105, square_with_reduction_special_prime_1_106, square_with_reduction_special_prime_1_107, square_with_reduction_special_prime_1_108, square_with_reduction_special_prime_1_109, square_with_reduction_special_prime_1_110, square_with_reduction_special_prime_1_111, square_with_reduction_special_prime_1_112, square_with_reduction_special_prime_1_113, square_with_reduction_special_prime_1_114, square_with_reduction_special_prime_1_115, square_with_reduction_special_prime_1_116, square_with_reduction_special_prime_1_117, square_with_reduction_special_prime_1_118, square_with_reduction_special_prime_1_119, square_with_reduction_special_prime_1_120, square_with_reduction_special_prime_1_121, square_with_reduction_special_prime_1_122, square_with_reduction_special_prime_1_123, square_with_reduction_special_prime_1_124, square_with_reduction_special_prime_1_125, square_with_reduction_special_prime_1_126, square_with_reduction_special_prime_1_127, square_with_reduction_special_prime_1_128, square_with_reduction_special_prime_1_129, square_with_reduction_special_prime_1_130, square_with_reduction_special_prime_1_131, square_with_reduction_special_prime_1_132, square_with_reduction_special_prime_1_133, square_with_reduction_special_prime_1_134, square_with_reduction_special_prime_1_135, square_with_reduction_special_prime_1_136, square_with_reduction_special_prime_1_137, square_with_reduction_special_prime_1_138, square_with_reduction_special_prime_1_139, 
square_with_reduction_special_prime_1_141, square_with_reduction_special_prime_1_142, square_with_reduction_special_prime_1_143, square_with_reduction_special_prime_1_144, square_with_reduction_special_prime_1_145, square_with_reduction_special_prime_1_146, square_with_reduction_special_prime_1_147, square_with_reduction_special_prime_1_148, square_with_reduction_special_prime_1_149, square_with_reduction_special_prime_1_150, square_with_reduction_special_prime_1_151, square_with_reduction_special_prime_1_152, square_with_reduction_special_prime_1_153, square_with_reduction_special_prime_1_154, square_with_reduction_special_prime_1_155, square_with_reduction_special_prime_1_156, square_with_reduction_special_prime_1_157, square_with_reduction_special_prime_1_158, square_with_reduction_special_prime_1_159, square_with_reduction_special_prime_1_160, square_with_reduction_special_prime_1_161, square_with_reduction_special_prime_1_162, square_with_reduction_special_prime_1_163, square_with_reduction_special_prime_1_164, square_with_reduction_special_prime_1_165, square_with_reduction_special_prime_1_166, square_with_reduction_special_prime_1_167, square_with_reduction_special_prime_1_168, square_with_reduction_special_prime_1_169, square_with_reduction_special_prime_1_170, square_with_reduction_special_prime_1_171, square_with_reduction_special_prime_1_172, square_with_reduction_special_prime_1_173, square_with_reduction_special_prime_1_174, square_with_reduction_special_prime_1_175, square_with_reduction_special_prime_1_176, square_with_reduction_special_prime_1_177, square_with_reduction_special_prime_1_178, square_with_reduction_special_prime_1_179, square_with_reduction_special_prime_1_180, square_with_reduction_special_prime_1_181, square_with_reduction_special_prime_1_182, square_with_reduction_special_prime_1_183, square_with_reduction_special_prime_1_184, square_with_reduction_special_prime_1_185, square_with_reduction_special_prime_1_186, square_with_reduction_special_prime_1_187, square_with_reduction_special_prime_1_188, square_with_reduction_special_prime_1_189, square_with_reduction_special_prime_1_190, square_with_reduction_special_prime_1_191, square_with_reduction_special_prime_1_192, square_with_reduction_special_prime_1_193, square_with_reduction_special_prime_1_194, square_with_reduction_special_prime_1_195, square_with_reduction_special_prime_1_196, 
square_with_reduction_special_prime_2_0, square_with_reduction_special_prime_2_1, square_with_reduction_special_prime_2_2, 
square_with_reduction_special_prime_2_4, square_with_reduction_special_prime_2_5, square_with_reduction_special_prime_2_6, square_with_reduction_special_prime_2_7, square_with_reduction_special_prime_2_8, square_with_reduction_special_prime_2_9, square_with_reduction_special_prime_2_10, square_with_reduction_special_prime_2_11, 
square_with_reduction_special_prime_2_13, square_with_reduction_special_prime_2_14, square_with_reduction_special_prime_2_15, square_with_reduction_special_prime_2_16, square_with_reduction_special_prime_2_17, square_with_reduction_special_prime_2_18, square_with_reduction_special_prime_2_19, square_with_reduction_special_prime_2_20, square_with_reduction_special_prime_2_21, square_with_reduction_special_prime_2_22, square_with_reduction_special_prime_2_23, square_with_reduction_special_prime_2_24, square_with_reduction_special_prime_2_25, square_with_reduction_special_prime_2_26, 
square_with_reduction_special_prime_2_28, square_with_reduction_special_prime_2_29, square_with_reduction_special_prime_2_30, square_with_reduction_special_prime_2_31, square_with_reduction_special_prime_2_32, square_with_reduction_special_prime_2_33, square_with_reduction_special_prime_2_34, square_with_reduction_special_prime_2_35, square_with_reduction_special_prime_2_36, square_with_reduction_special_prime_2_37, square_with_reduction_special_prime_2_38, square_with_reduction_special_prime_2_39, square_with_reduction_special_prime_2_40, square_with_reduction_special_prime_2_41, square_with_reduction_special_prime_2_42, square_with_reduction_special_prime_2_43, square_with_reduction_special_prime_2_44, square_with_reduction_special_prime_2_45, square_with_reduction_special_prime_2_46, square_with_reduction_special_prime_2_47, square_with_reduction_special_prime_2_48, square_with_reduction_special_prime_2_49,
square_with_reduction_special_prime_2_51, square_with_reduction_special_prime_2_52, square_with_reduction_special_prime_2_53, square_with_reduction_special_prime_2_54, square_with_reduction_special_prime_2_55, square_with_reduction_special_prime_2_56, square_with_reduction_special_prime_2_57, square_with_reduction_special_prime_2_58, square_with_reduction_special_prime_2_59, square_with_reduction_special_prime_2_60, square_with_reduction_special_prime_2_61, square_with_reduction_special_prime_2_62, square_with_reduction_special_prime_2_63, square_with_reduction_special_prime_2_64, square_with_reduction_special_prime_2_65, square_with_reduction_special_prime_2_66, square_with_reduction_special_prime_2_67, square_with_reduction_special_prime_2_68, square_with_reduction_special_prime_2_69, square_with_reduction_special_prime_2_70, square_with_reduction_special_prime_2_71, square_with_reduction_special_prime_2_72, square_with_reduction_special_prime_2_73, square_with_reduction_special_prime_2_74, square_with_reduction_special_prime_2_75, square_with_reduction_special_prime_2_76, square_with_reduction_special_prime_2_77, square_with_reduction_special_prime_2_78, square_with_reduction_special_prime_2_79, square_with_reduction_special_prime_2_80, square_with_reduction_special_prime_2_81,
square_with_reduction_special_prime_2_83, square_with_reduction_special_prime_2_84, square_with_reduction_special_prime_2_85, square_with_reduction_special_prime_2_86, square_with_reduction_special_prime_2_87, square_with_reduction_special_prime_2_88, square_with_reduction_special_prime_2_89, square_with_reduction_special_prime_2_90, square_with_reduction_special_prime_2_91, square_with_reduction_special_prime_2_92, square_with_reduction_special_prime_2_93, square_with_reduction_special_prime_2_94, square_with_reduction_special_prime_2_95, square_with_reduction_special_prime_2_96, square_with_reduction_special_prime_2_97, square_with_reduction_special_prime_2_98, square_with_reduction_special_prime_2_99, square_with_reduction_special_prime_2_100, square_with_reduction_special_prime_2_101, square_with_reduction_special_prime_2_102, square_with_reduction_special_prime_2_103, square_with_reduction_special_prime_2_104, square_with_reduction_special_prime_2_105, square_with_reduction_special_prime_2_106, square_with_reduction_special_prime_2_107, square_with_reduction_special_prime_2_108, square_with_reduction_special_prime_2_109, square_with_reduction_special_prime_2_110, square_with_reduction_special_prime_2_111, square_with_reduction_special_prime_2_112, square_with_reduction_special_prime_2_113, square_with_reduction_special_prime_2_114, square_with_reduction_special_prime_2_115, square_with_reduction_special_prime_2_116, square_with_reduction_special_prime_2_117, square_with_reduction_special_prime_2_118, square_with_reduction_special_prime_2_119, square_with_reduction_special_prime_2_120, square_with_reduction_special_prime_2_121, square_with_reduction_special_prime_2_122, square_with_reduction_special_prime_2_123, square_with_reduction_special_prime_2_124, 
 square_with_reduction_special_prime_2_126, square_with_reduction_special_prime_2_127, square_with_reduction_special_prime_2_128, square_with_reduction_special_prime_2_129, square_with_reduction_special_prime_2_130, square_with_reduction_special_prime_2_131, square_with_reduction_special_prime_2_132, square_with_reduction_special_prime_2_133, square_with_reduction_special_prime_2_134, square_with_reduction_special_prime_2_135, square_with_reduction_special_prime_2_136, square_with_reduction_special_prime_2_137, square_with_reduction_special_prime_2_138, square_with_reduction_special_prime_2_139, square_with_reduction_special_prime_2_140, square_with_reduction_special_prime_2_141, square_with_reduction_special_prime_2_142, square_with_reduction_special_prime_2_143, square_with_reduction_special_prime_2_144, square_with_reduction_special_prime_2_145, square_with_reduction_special_prime_2_146, square_with_reduction_special_prime_2_147, square_with_reduction_special_prime_2_148, square_with_reduction_special_prime_2_149, square_with_reduction_special_prime_2_150, square_with_reduction_special_prime_2_151, square_with_reduction_special_prime_2_152, square_with_reduction_special_prime_2_153, square_with_reduction_special_prime_2_154, square_with_reduction_special_prime_2_155, square_with_reduction_special_prime_2_156, square_with_reduction_special_prime_2_157, square_with_reduction_special_prime_2_158, square_with_reduction_special_prime_2_159, square_with_reduction_special_prime_2_160, square_with_reduction_special_prime_2_161, square_with_reduction_special_prime_2_162, square_with_reduction_special_prime_2_163, square_with_reduction_special_prime_2_164, square_with_reduction_special_prime_2_165, square_with_reduction_special_prime_2_166, square_with_reduction_special_prime_2_167, square_with_reduction_special_prime_2_168, square_with_reduction_special_prime_2_169, square_with_reduction_special_prime_2_170, square_with_reduction_special_prime_2_171, square_with_reduction_special_prime_2_172, square_with_reduction_special_prime_2_173, square_with_reduction_special_prime_2_174, square_with_reduction_special_prime_2_175, square_with_reduction_special_prime_2_176, square_with_reduction_special_prime_2_177, square_with_reduction_special_prime_2_178, square_with_reduction_special_prime_2_179, 
square_with_reduction_special_prime_3_0, square_with_reduction_special_prime_3_1, square_with_reduction_special_prime_3_2, square_with_reduction_special_prime_3_3, square_with_reduction_special_prime_3_4, square_with_reduction_special_prime_3_5, 
square_with_reduction_special_prime_3_7, square_with_reduction_special_prime_3_8, square_with_reduction_special_prime_3_9, square_with_reduction_special_prime_3_10, square_with_reduction_special_prime_3_11, square_with_reduction_special_prime_3_12, square_with_reduction_special_prime_3_13, square_with_reduction_special_prime_3_14, square_with_reduction_special_prime_3_15, square_with_reduction_special_prime_3_16, square_with_reduction_special_prime_3_17, 
square_with_reduction_special_prime_3_19, square_with_reduction_special_prime_3_20, square_with_reduction_special_prime_3_21, square_with_reduction_special_prime_3_22, square_with_reduction_special_prime_3_23, square_with_reduction_special_prime_3_24, square_with_reduction_special_prime_3_25, square_with_reduction_special_prime_3_26, square_with_reduction_special_prime_3_27, square_with_reduction_special_prime_3_28, square_with_reduction_special_prime_3_29, square_with_reduction_special_prime_3_30, square_with_reduction_special_prime_3_31, square_with_reduction_special_prime_3_32, square_with_reduction_special_prime_3_33, square_with_reduction_special_prime_3_34, square_with_reduction_special_prime_3_35, square_with_reduction_special_prime_3_36, square_with_reduction_special_prime_3_37, 
square_with_reduction_special_prime_3_39, square_with_reduction_special_prime_3_40, square_with_reduction_special_prime_3_41, square_with_reduction_special_prime_3_42, square_with_reduction_special_prime_3_43, square_with_reduction_special_prime_3_44, square_with_reduction_special_prime_3_45, square_with_reduction_special_prime_3_46, square_with_reduction_special_prime_3_47, square_with_reduction_special_prime_3_48, square_with_reduction_special_prime_3_49, square_with_reduction_special_prime_3_50, square_with_reduction_special_prime_3_51, square_with_reduction_special_prime_3_52, square_with_reduction_special_prime_3_53, square_with_reduction_special_prime_3_54, square_with_reduction_special_prime_3_55, square_with_reduction_special_prime_3_56, square_with_reduction_special_prime_3_57, square_with_reduction_special_prime_3_58, square_with_reduction_special_prime_3_59, square_with_reduction_special_prime_3_60, square_with_reduction_special_prime_3_61, square_with_reduction_special_prime_3_62, square_with_reduction_special_prime_3_63, square_with_reduction_special_prime_3_64, square_with_reduction_special_prime_3_65, square_with_reduction_special_prime_3_66, 
square_with_reduction_special_prime_3_68, square_with_reduction_special_prime_3_69, square_with_reduction_special_prime_3_70, square_with_reduction_special_prime_3_71, square_with_reduction_special_prime_3_72, square_with_reduction_special_prime_3_73, square_with_reduction_special_prime_3_74, square_with_reduction_special_prime_3_75, square_with_reduction_special_prime_3_76, square_with_reduction_special_prime_3_77, square_with_reduction_special_prime_3_78, square_with_reduction_special_prime_3_79, square_with_reduction_special_prime_3_80, square_with_reduction_special_prime_3_81, square_with_reduction_special_prime_3_82, square_with_reduction_special_prime_3_83, square_with_reduction_special_prime_3_84, square_with_reduction_special_prime_3_85, square_with_reduction_special_prime_3_86, square_with_reduction_special_prime_3_87, square_with_reduction_special_prime_3_88, square_with_reduction_special_prime_3_89, square_with_reduction_special_prime_3_90, square_with_reduction_special_prime_3_91, square_with_reduction_special_prime_3_92, square_with_reduction_special_prime_3_93, square_with_reduction_special_prime_3_94, square_with_reduction_special_prime_3_95, square_with_reduction_special_prime_3_96, square_with_reduction_special_prime_3_97, square_with_reduction_special_prime_3_98, square_with_reduction_special_prime_3_99, square_with_reduction_special_prime_3_100, square_with_reduction_special_prime_3_101, square_with_reduction_special_prime_3_102, square_with_reduction_special_prime_3_103, square_with_reduction_special_prime_3_104, square_with_reduction_special_prime_3_105, square_with_reduction_special_prime_3_106,
square_with_reduction_special_prime_3_108, square_with_reduction_special_prime_3_109, square_with_reduction_special_prime_3_110, square_with_reduction_special_prime_3_111, square_with_reduction_special_prime_3_112, square_with_reduction_special_prime_3_113, square_with_reduction_special_prime_3_114, square_with_reduction_special_prime_3_115, square_with_reduction_special_prime_3_116, square_with_reduction_special_prime_3_117, square_with_reduction_special_prime_3_118, square_with_reduction_special_prime_3_119, square_with_reduction_special_prime_3_120, square_with_reduction_special_prime_3_121, square_with_reduction_special_prime_3_122, square_with_reduction_special_prime_3_123, square_with_reduction_special_prime_3_124, square_with_reduction_special_prime_3_125, square_with_reduction_special_prime_3_126, square_with_reduction_special_prime_3_127, square_with_reduction_special_prime_3_128, square_with_reduction_special_prime_3_129, square_with_reduction_special_prime_3_130, square_with_reduction_special_prime_3_131, square_with_reduction_special_prime_3_132, square_with_reduction_special_prime_3_133, square_with_reduction_special_prime_3_134, square_with_reduction_special_prime_3_135, square_with_reduction_special_prime_3_136, square_with_reduction_special_prime_3_137, square_with_reduction_special_prime_3_138, square_with_reduction_special_prime_3_139, square_with_reduction_special_prime_3_140, square_with_reduction_special_prime_3_141, square_with_reduction_special_prime_3_142, square_with_reduction_special_prime_3_143, square_with_reduction_special_prime_3_144, square_with_reduction_special_prime_3_145, square_with_reduction_special_prime_3_146, square_with_reduction_special_prime_3_147, square_with_reduction_special_prime_3_148, square_with_reduction_special_prime_3_149, square_with_reduction_special_prime_3_150, square_with_reduction_special_prime_3_151, square_with_reduction_special_prime_3_152, square_with_reduction_special_prime_3_153, square_with_reduction_special_prime_3_154, square_with_reduction_special_prime_3_155, square_with_reduction_special_prime_3_156, square_with_reduction_special_prime_3_157, square_with_reduction_special_prime_3_158,
-- 0100 addition/subtraction with no reduction
addition_subtraction_direct_0, addition_subtraction_direct_2, addition_subtraction_direct_3, addition_subtraction_direct_5, addition_subtraction_direct_6, addition_subtraction_direct_8, addition_subtraction_direct_9, addition_subtraction_direct_11, addition_subtraction_direct_12, addition_subtraction_direct_14, addition_subtraction_direct_15, addition_subtraction_direct_17, addition_subtraction_direct_18, addition_subtraction_direct_20, addition_subtraction_direct_21,
-- 0101 iterative modular reduction
iterative_modular_reduction_0, iterative_modular_reduction_1, iterative_modular_reduction_2, iterative_modular_reduction_3,
iterative_modular_reduction_5, iterative_modular_reduction_6, iterative_modular_reduction_7, iterative_modular_reduction_8, iterative_modular_reduction_9, iterative_modular_reduction_10, iterative_modular_reduction_11,
iterative_modular_reduction_13, iterative_modular_reduction_14, iterative_modular_reduction_15, iterative_modular_reduction_16, iterative_modular_reduction_17, iterative_modular_reduction_18, iterative_modular_reduction_19, iterative_modular_reduction_20, iterative_modular_reduction_21, iterative_modular_reduction_22,
iterative_modular_reduction_24, iterative_modular_reduction_25, iterative_modular_reduction_26, iterative_modular_reduction_27, iterative_modular_reduction_28, iterative_modular_reduction_29, iterative_modular_reduction_30, iterative_modular_reduction_31, iterative_modular_reduction_32, iterative_modular_reduction_33, iterative_modular_reduction_34, iterative_modular_reduction_35, iterative_modular_reduction_36,
iterative_modular_reduction_38, iterative_modular_reduction_39, iterative_modular_reduction_40, iterative_modular_reduction_41, iterative_modular_reduction_42, iterative_modular_reduction_43, iterative_modular_reduction_44, iterative_modular_reduction_45, iterative_modular_reduction_46, iterative_modular_reduction_47, iterative_modular_reduction_48, iterative_modular_reduction_49, iterative_modular_reduction_50, iterative_modular_reduction_51, iterative_modular_reduction_52, iterative_modular_reduction_53,
iterative_modular_reduction_55, iterative_modular_reduction_56, iterative_modular_reduction_57, iterative_modular_reduction_58, iterative_modular_reduction_59, iterative_modular_reduction_60, iterative_modular_reduction_61, iterative_modular_reduction_62, iterative_modular_reduction_63, iterative_modular_reduction_64, iterative_modular_reduction_65, iterative_modular_reduction_66, iterative_modular_reduction_67, iterative_modular_reduction_68, iterative_modular_reduction_69, iterative_modular_reduction_70, iterative_modular_reduction_71, iterative_modular_reduction_72, iterative_modular_reduction_73,
iterative_modular_reduction_75, iterative_modular_reduction_76, iterative_modular_reduction_77, iterative_modular_reduction_78, iterative_modular_reduction_79, iterative_modular_reduction_80, iterative_modular_reduction_81, iterative_modular_reduction_82, iterative_modular_reduction_83, iterative_modular_reduction_84, iterative_modular_reduction_85, iterative_modular_reduction_86, iterative_modular_reduction_87, iterative_modular_reduction_88, iterative_modular_reduction_89, iterative_modular_reduction_90, iterative_modular_reduction_91, iterative_modular_reduction_92, iterative_modular_reduction_93, iterative_modular_reduction_94, iterative_modular_reduction_95, iterative_modular_reduction_96,
iterative_modular_reduction_98, iterative_modular_reduction_99, iterative_modular_reduction_100, iterative_modular_reduction_101, iterative_modular_reduction_102, iterative_modular_reduction_103, iterative_modular_reduction_104, iterative_modular_reduction_105, iterative_modular_reduction_106, iterative_modular_reduction_107, iterative_modular_reduction_108, iterative_modular_reduction_109, iterative_modular_reduction_110, iterative_modular_reduction_111, iterative_modular_reduction_112, iterative_modular_reduction_113, iterative_modular_reduction_114, iterative_modular_reduction_115, iterative_modular_reduction_116, iterative_modular_reduction_117, iterative_modular_reduction_118, iterative_modular_reduction_119, iterative_modular_reduction_120, iterative_modular_reduction_121, iterative_modular_reduction_122,
-- 0110 addition/subtraction with reduction
addition_subtraction_with_reduction_0, addition_subtraction_with_reduction_1, addition_subtraction_with_reduction_2, addition_subtraction_with_reduction_3,
addition_subtraction_with_reduction_5, addition_subtraction_with_reduction_6, addition_subtraction_with_reduction_7, addition_subtraction_with_reduction_8, addition_subtraction_with_reduction_9, addition_subtraction_with_reduction_10, addition_subtraction_with_reduction_11, addition_subtraction_with_reduction_12,
addition_subtraction_with_reduction_14, addition_subtraction_with_reduction_15, addition_subtraction_with_reduction_16, addition_subtraction_with_reduction_17, addition_subtraction_with_reduction_18, addition_subtraction_with_reduction_19, addition_subtraction_with_reduction_20, addition_subtraction_with_reduction_21, addition_subtraction_with_reduction_22, addition_subtraction_with_reduction_23, addition_subtraction_with_reduction_24,
addition_subtraction_with_reduction_26, addition_subtraction_with_reduction_27, addition_subtraction_with_reduction_28, addition_subtraction_with_reduction_29, addition_subtraction_with_reduction_30, addition_subtraction_with_reduction_31, addition_subtraction_with_reduction_32, addition_subtraction_with_reduction_33, addition_subtraction_with_reduction_34, addition_subtraction_with_reduction_35, addition_subtraction_with_reduction_36, addition_subtraction_with_reduction_37, addition_subtraction_with_reduction_38, addition_subtraction_with_reduction_39,
addition_subtraction_with_reduction_41, addition_subtraction_with_reduction_42, addition_subtraction_with_reduction_43, addition_subtraction_with_reduction_44, addition_subtraction_with_reduction_45, addition_subtraction_with_reduction_46, addition_subtraction_with_reduction_47, addition_subtraction_with_reduction_48, addition_subtraction_with_reduction_49, addition_subtraction_with_reduction_50, addition_subtraction_with_reduction_51, addition_subtraction_with_reduction_52, addition_subtraction_with_reduction_53, addition_subtraction_with_reduction_54, addition_subtraction_with_reduction_55, addition_subtraction_with_reduction_56, addition_subtraction_with_reduction_57,
addition_subtraction_with_reduction_59, addition_subtraction_with_reduction_60, addition_subtraction_with_reduction_61, addition_subtraction_with_reduction_62, addition_subtraction_with_reduction_63, addition_subtraction_with_reduction_64, addition_subtraction_with_reduction_65, addition_subtraction_with_reduction_66, addition_subtraction_with_reduction_67, addition_subtraction_with_reduction_68, addition_subtraction_with_reduction_69, addition_subtraction_with_reduction_70, addition_subtraction_with_reduction_71, addition_subtraction_with_reduction_72, addition_subtraction_with_reduction_73, addition_subtraction_with_reduction_74, addition_subtraction_with_reduction_75, addition_subtraction_with_reduction_76, addition_subtraction_with_reduction_77, addition_subtraction_with_reduction_78,
addition_subtraction_with_reduction_80, addition_subtraction_with_reduction_81, addition_subtraction_with_reduction_82, addition_subtraction_with_reduction_83, addition_subtraction_with_reduction_84, addition_subtraction_with_reduction_85, addition_subtraction_with_reduction_86, addition_subtraction_with_reduction_87, addition_subtraction_with_reduction_88, addition_subtraction_with_reduction_89, addition_subtraction_with_reduction_90, addition_subtraction_with_reduction_91, addition_subtraction_with_reduction_92, addition_subtraction_with_reduction_93, addition_subtraction_with_reduction_94, addition_subtraction_with_reduction_95, addition_subtraction_with_reduction_96, addition_subtraction_with_reduction_97, addition_subtraction_with_reduction_98, addition_subtraction_with_reduction_99, addition_subtraction_with_reduction_100, addition_subtraction_with_reduction_101, addition_subtraction_with_reduction_102,
addition_subtraction_with_reduction_104, addition_subtraction_with_reduction_105, addition_subtraction_with_reduction_106, addition_subtraction_with_reduction_107, addition_subtraction_with_reduction_108, addition_subtraction_with_reduction_109, addition_subtraction_with_reduction_110, addition_subtraction_with_reduction_111, addition_subtraction_with_reduction_112, addition_subtraction_with_reduction_113, addition_subtraction_with_reduction_114, addition_subtraction_with_reduction_115, addition_subtraction_with_reduction_116, addition_subtraction_with_reduction_117, addition_subtraction_with_reduction_118, addition_subtraction_with_reduction_119, addition_subtraction_with_reduction_120, addition_subtraction_with_reduction_121, addition_subtraction_with_reduction_122, addition_subtraction_with_reduction_123, addition_subtraction_with_reduction_124, addition_subtraction_with_reduction_125, addition_subtraction_with_reduction_126, addition_subtraction_with_reduction_127, addition_subtraction_with_reduction_128, addition_subtraction_with_reduction_129,
-- NOP
nop_4_stages, nop_8_stages
); 

signal actual_state, next_state : state;

signal next_sm_rotation_size : std_logic_vector(1 downto 0);
signal next_sm_circular_shift_enable : std_logic;
signal next_sel_address_a : std_logic;
signal next_sel_address_b_prime : std_logic_vector(1 downto 0);
signal next_sm_specific_mac_address_a : std_logic_vector(2 downto 0);
signal next_sm_specific_mac_address_b : std_logic_vector(2 downto 0);
signal next_sm_specific_mac_address_o : std_logic_vector(2 downto 0);
signal next_sm_specific_mac_next_address_o : std_logic_vector(2 downto 0);
signal next_mac_enable_signed_a : std_logic;
signal next_mac_enable_signed_b : std_logic;
signal next_mac_sel_load_reg_a : std_logic_vector(1 downto 0);
signal next_mac_clear_reg_b : std_logic;
signal next_mac_clear_reg_acc : std_logic;
signal next_mac_sel_shift_reg_o : std_logic;
signal next_mac_enable_update_reg_s : std_logic;
signal next_mac_sel_reg_s_reg_o_sign : std_logic;
signal next_mac_reg_s_reg_o_positive : std_logic;
signal next_sm_sign_a_mode : std_logic;
signal next_sm_mac_operation_mode : std_logic_vector(1 downto 0);
signal next_mac_enable_reg_s_mask : std_logic;
signal next_mac_subtraction_reg_a_b : std_logic;
signal next_mac_sel_multiply_two_a_b : std_logic;
signal next_mac_sel_reg_y_output : std_logic;
signal next_sm_mac_write_enable_output : std_logic;
signal next_mac_memory_double_mode : std_logic;
signal next_mac_memory_only_write_mode : std_logic;
signal next_base_address_generator_o_increment_previous_address : std_logic;
signal next_sm_free_flag : std_logic;

signal ultimate_operation : std_logic;

begin

process(clk)
begin
    if(rising_edge(clk)) then
        if(rstn = '0') then
            ultimate_operation <= '0';
        else
            ultimate_operation <= penultimate_operation;
        end if;
    end if;
end process;

registers_state : process(clk, rstn)
begin
    if(rstn = '0') then
        actual_state <= reset;
    elsif(rising_edge(clk)) then
        actual_state <= next_state;
    end if;
end process;

registers_state_output : process(clk)
begin
    if(rising_edge(clk)) then
        if(rstn = '0') then
            sm_free_flag <= '0';
            sm_rotation_size <= "11";
            sm_circular_shift_enable <= '0';
            sel_address_a <= '0';
            sel_address_b_prime <= "00";
            sm_specific_mac_address_a <= "000";
            sm_specific_mac_address_b <= "000";
            sm_specific_mac_address_o <= "000";
            sm_specific_mac_next_address_o <= "001";
            mac_enable_signed_a <= '0';
            mac_enable_signed_b <= '0';
            mac_sel_load_reg_a <= "11";
            mac_clear_reg_b <= '1';
            mac_clear_reg_acc <= '1';
            mac_sel_shift_reg_o <= '0';
            mac_enable_update_reg_s <= '0';
            mac_sel_reg_s_reg_o_sign <= '0';
            mac_reg_s_reg_o_positive <= '0';
            sm_sign_a_mode <= '0';
            sm_mac_operation_mode <= "10";
            mac_enable_reg_s_mask <= '0';
            mac_subtraction_reg_a_b <= '0';
            mac_sel_multiply_two_a_b <= '0';
            mac_sel_reg_y_output <= '0';
            base_address_generator_o_increment_previous_address <= '0';
            sm_mac_write_enable_output <= '0';
            mac_memory_double_mode <= '0';
            mac_memory_only_write_mode <= '0';
        else
            sm_free_flag <= next_sm_free_flag;
            sm_rotation_size <= next_sm_rotation_size;
            sm_circular_shift_enable <= next_sm_circular_shift_enable;
            sel_address_a <= next_sel_address_a;
            sel_address_b_prime <= next_sel_address_b_prime;
            sm_specific_mac_address_a <= next_sm_specific_mac_address_a;
            sm_specific_mac_address_b <= next_sm_specific_mac_address_b;
            sm_specific_mac_address_o <= next_sm_specific_mac_address_o;
            sm_specific_mac_next_address_o <= next_sm_specific_mac_next_address_o;
            mac_enable_signed_a <= next_mac_enable_signed_a;
            mac_enable_signed_b <= next_mac_enable_signed_b;
            mac_sel_load_reg_a <= next_mac_sel_load_reg_a;
            mac_clear_reg_b <= next_mac_clear_reg_b;
            mac_clear_reg_acc <= next_mac_clear_reg_acc;
            mac_sel_shift_reg_o <= next_mac_sel_shift_reg_o;
            mac_enable_update_reg_s <= next_mac_enable_update_reg_s;
            mac_sel_reg_s_reg_o_sign <= next_mac_sel_reg_s_reg_o_sign;
            mac_reg_s_reg_o_positive <= next_mac_reg_s_reg_o_positive;
            sm_sign_a_mode <= next_sm_sign_a_mode;
            sm_mac_operation_mode <= next_sm_mac_operation_mode;
            mac_enable_reg_s_mask <= next_mac_enable_reg_s_mask;
            mac_subtraction_reg_a_b <= next_mac_subtraction_reg_a_b;
            mac_sel_multiply_two_a_b <= next_mac_sel_multiply_two_a_b;
            mac_sel_reg_y_output <= next_mac_sel_reg_y_output;
            base_address_generator_o_increment_previous_address <= next_base_address_generator_o_increment_previous_address;
            sm_mac_write_enable_output <= next_sm_mac_write_enable_output;
            mac_memory_double_mode <= next_mac_memory_double_mode;
            mac_memory_only_write_mode <= next_mac_memory_only_write_mode;
        end if;
    end if;
end process;

update_output : process(next_state)
begin
    case (next_state) is
        when reset =>
            next_sm_free_flag <= '1';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '0';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "11";
            next_mac_clear_reg_b <= '1';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when decode_instruction =>
            next_sm_free_flag <= '1';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '0';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "11";
            next_mac_clear_reg_b <= '1';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_0 =>
            -- -- In case of size 1
            -- reg_a = a0_X; reg_b = b0_X; reg_acc = 0; o0_X = reg_o; o1_X = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_2 =>
            -- -- Other cases
            -- reg_a = a0_X; reg_b = b0_X; reg_acc = 0; o0_X = reg_o; operation : a*b + acc; o0_X = reg_o;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_3 =>
            -- -- In case of size 2
            -- reg_a = a1_X; reg_b = b0_X; reg_acc = reg_o >> 256; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_4 =>
            -- reg_a = a0_X; reg_b = b1_X; reg_acc = reg_o; o1_X = reg_o; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_5 =>
            -- reg_a = a1_X; reg_b = b1_X; reg_acc = reg_o >> 256; o2_X = reg_o; o3_X = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_7 =>
            -- -- Other cases
            -- reg_a = a1_X; reg_b = b0_X; reg_acc = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_8 =>
            -- reg_a = a0_X; reg_b = b1_X; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_9 =>
            -- reg_a = a1_X; reg_b = b1_X; reg_acc = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_10 =>
            -- -- In case of size 3
            -- reg_a = a0_X; reg_b = b2_X; reg_acc = reg_o; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_11 =>
            -- reg_a = a2_X; reg_b = b0_X; reg_acc = reg_o; Enable sign a; o2_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_12 =>
            -- reg_a = a2_X; reg_b = b1_X; reg_acc = reg_o >> 256; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_13 =>
            -- reg_a = a1_X; reg_b = b2_X; reg_acc = reg_o; o3_X = reg_o; Enable sign b; operation : a*b + acc; 
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_14 =>
            -- reg_a = a2_X; reg_b = b2_X; reg_acc = reg_o >> 256; o4_X = reg_o; o5_X = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_16 =>
            -- -- Other cases
            -- reg_a = a0_0; reg_b = b2_0; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_17 =>
            -- reg_a = a2_X; reg_b = b0_X; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_18 =>
            -- reg_a = a2_X; reg_b = b1_X; reg_acc = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_19 =>
            -- reg_a = a1_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc; 
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_20 =>
            -- -- In case of size 4
            -- reg_a = a3_X; reg_b = b0_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_21 =>
            -- reg_a = a0_X; reg_b = b3_X; reg_acc = reg_o; o3_X = reg_o; Enable sign b; operation : a*b + acc; 
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_22 =>
            -- reg_a = a2_X; reg_b = b2_X; reg_acc = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_23 =>
            -- reg_a = a3_X; reg_b = b1_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_24 =>
            -- reg_a = a1_X; reg_b = b3_X; reg_acc = reg_o; o4_X = reg_o; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_25 =>
            -- reg_a = a3_X; reg_b = b2_X; reg_acc = reg_o >> 256; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_26 =>
            -- reg_a = a2_X; reg_b = b3_X; reg_acc = reg_o; o5_X = reg_o; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_27 =>
            -- reg_a = a3_X; reg_b = b3_X; reg_acc = reg_o >> 256; o6_X = reg_o; o7_X = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_29 =>
            -- -- Other cases
            -- reg_a = a3_X; reg_b = b0_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_30 =>
            -- reg_a = a0_X; reg_b = b3_X; reg_acc = reg_o; o3_0 = reg_o; operation : a*b + acc; 
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_31 =>
            -- reg_a = a2_X; reg_b = b2_X; reg_acc = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_32 =>
            -- reg_a = a3_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_33 =>
            -- reg_a = a1_X; reg_b = b3_X; reg_acc = reg_o; o4_0 = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_34 =>
            -- -- In case of size 5
            -- reg_a = a4_X; reg_b = b0_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_35 =>
            -- reg_a = a0_X; reg_b = b4_X; reg_acc = reg_o; o4_0 = reg_o; Enable sign b; operation : a*b + acc; 
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_36 =>
            -- reg_a = a3_X; reg_b = b2_X; reg_acc = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_37 =>
            -- reg_a = a2_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_38 =>
            -- reg_a = a4_X; reg_b = b1_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_39 =>
            -- reg_a = a1_X; reg_b = b4_X; reg_acc = reg_o; o5_X = reg_o; Enable sign b; operation : a*b + acc; 
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_40 =>
            -- reg_a = a3_X; reg_b = b3_X; reg_acc = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_41 =>
            -- reg_a = a4_X; reg_b = b2_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_42 =>
            -- reg_a = a2_X; reg_b = b4_X; reg_acc = reg_o; o6_X = reg_o; Enable sign b; operation : a*b + acc; 
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_43 =>
            -- reg_a = a4_X; reg_b = b3_X; reg_acc = reg_o >> 256; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "111";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_44 =>
            -- reg_a = a3_X; reg_b = b4_X; reg_acc = reg_o; o7_X = reg_o; Enable sign b; operation : a*b + acc; Increment base address o;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "111";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '1';
        when multiplication_direct_45 =>
            -- reg_a = a4_X; reg_b = b4_X; reg_acc = reg_o >> 256; o8_X = reg_o; o9_X = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_47 =>
            -- -- Other cases
            -- reg_a = a4_X; reg_b = b0_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_48 =>
            -- reg_a = a0_X; reg_b = b4_X; reg_acc = reg_o; o4_X = reg_o; operation : a*b + acc; 
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_49 =>
            -- reg_a = a3_X; reg_b = b2_X; reg_acc = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_50 =>
            -- reg_a = a2_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_51 =>
            -- reg_a = a4_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_52 =>
            -- reg_a = a1_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc; 
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_53 =>
            -- -- In case of size 6
            -- reg_a = a5_X; reg_b = b0_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_54 =>
            -- reg_a = a0_X; reg_b = b5_X; reg_acc = reg_o; o5_0 = reg_o; Enable sign b; operation : a*b + acc; 
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_55 =>
            -- reg_a = a3_X; reg_b = b3_X; reg_acc = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_56 =>
            -- reg_a = a2_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_57 =>
            -- reg_a = a4_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_58 =>
            -- reg_a = a5_X; reg_b = b1_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_59 =>
            -- reg_a = a1_X; reg_b = b5_X; reg_acc = reg_o; o6_0 = reg_o; Enable sign b; operation : a*b + acc; 
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_60 =>
            -- reg_a = a4_X; reg_b = b3_X; reg_acc = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "111";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_61 =>
            -- reg_a = a3_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "111";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_62 =>
            -- reg_a = a5_X; reg_b = b2_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "111";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_63 =>
            -- reg_a = a2_X; reg_b = b5_X; reg_acc = reg_o; o7_0 = reg_o; Enable sign b; operation : a*b + acc; Increment base address o;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "111";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '1';
        when multiplication_direct_64 =>
            -- reg_a = a4_X; reg_b = b4_X; reg_acc = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_65 =>
            -- reg_a = a5_X; reg_b = b3_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_66 =>
            -- reg_a = a3_X; reg_b = b5_X; reg_acc = reg_o; o8_0 = reg_o; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_67 =>
            -- reg_a = a5_X; reg_b = b4_X; reg_acc = reg_o >> 256; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_68 =>
            -- reg_a = a4_X; reg_b = b5_X; reg_acc = reg_o; o9_0 = reg_o; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_69 =>
            -- reg_a = a5_X; reg_b = b5_X; reg_acc = reg_o >> 256; o10_X = reg_o; o11_X = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_71 =>
            -- -- Other cases
            -- reg_a = a5_X; reg_b = b0_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_72 =>
            -- reg_a = a0_X; reg_b = b5_X; reg_acc = reg_o; o5_0 = reg_o; operation : a*b + acc; 
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_73 =>
            -- reg_a = a3_X; reg_b = b3_X; reg_acc = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_74 =>
            -- reg_a = a4_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_75 =>
            -- reg_a = a2_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_76 =>
            -- reg_a = a5_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_77 =>
            -- reg_a = a1_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_78 =>
            -- -- In case of size 7
            -- reg_a = a6_X; reg_b = b0_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_79 =>
            -- reg_a = a0_X; reg_b = b6_X; reg_acc = reg_o; o6_0 = reg_o; Enable sign b; operation : a*b + acc; 
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_80 =>
            -- reg_a = a4_X; reg_b = b3_X; reg_acc = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "111";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_81 =>
            -- reg_a = a3_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "111";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_82 =>
            -- reg_a = a5_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "111";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_83 =>
            -- reg_a = a2_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "111";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_84 =>
            -- reg_a = a6_X; reg_b = b1_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "111";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_85 =>
            -- reg_a = a1_X; reg_b = b6_X; reg_acc = reg_o; o7_0 = reg_o; Enable sign b; operation : a*b + acc; Increment base address o;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "111";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '1';
        when multiplication_direct_86 =>
            -- reg_a = a4_X; reg_b = b4_X; reg_acc = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_87 =>
            -- reg_a = a5_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_88 =>
            -- reg_a = a3_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_89 =>
            -- reg_a = a6_X; reg_b = b2_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_90 =>
            -- reg_a = a2_X; reg_b = b6_X; reg_acc = reg_o; o8_0 = reg_o; Enable sign b; operation : a*b + acc; 
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_91 =>
            -- reg_a = a5_X; reg_b = b4_X; reg_acc = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_92 =>
            -- reg_a = a4_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_93 =>
            -- reg_a = a6_X; reg_b = b3_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_94 =>
            -- reg_a = a3_X; reg_b = b6_X; reg_acc = reg_o; o9_0 = reg_o; Enable sign b; operation : a*b + acc; 
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_95 =>
            -- reg_a = a5_X; reg_b = b5_X; reg_acc = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_96 =>
            -- reg_a = a6_X; reg_b = b4_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_97 =>
            -- reg_a = a4_X; reg_b = b6_X; reg_acc = reg_o; o10_0 = reg_o; Enable sign b; operation : a*b + acc; 
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_98 =>
            -- reg_a = a6_X; reg_b = b5_X; reg_acc = reg_o >> 256; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_99 =>
            -- reg_a = a5_X; reg_b = b6_X; reg_acc = reg_o; o11_0 = reg_o; Enable sign b; operation : a*b + acc; 
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_100 =>
            -- reg_a = a6_X; reg_b = b6_X; reg_acc = reg_o >> 256; o12_X = reg_o; o13_X = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_102 =>
            -- -- In case of size 8
            -- reg_a = a6_X; reg_b = b0_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_103 =>
            -- reg_a = a0_X; reg_b = b6_X; reg_acc = reg_o; o6_0 = reg_o; operation : a*b + acc; 
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_104 =>
            -- reg_a = a4_X; reg_b = b3_X; reg_acc = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "111";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_105 =>
            -- reg_a = a3_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "111";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_106 =>
            -- reg_a = a5_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "111";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_107 =>
            -- reg_a = a2_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "111";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_108 =>
            -- reg_a = a6_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "111";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_109 =>
            -- reg_a = a1_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "111";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_110 =>
            -- reg_a = a7_X; reg_b = b0_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "111";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_111 =>
            -- reg_a = a0_X; reg_b = b7_X; reg_acc = reg_o; o7_0 = reg_o; Enable sign b; operation : a*b + acc; Increment base address o;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "111";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '1';
        when multiplication_direct_112 =>
            -- reg_a = a4_X; reg_b = b4_X; reg_acc = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_113 =>
            -- reg_a = a5_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_114 =>
            -- reg_a = a3_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_115 =>
            -- reg_a = a6_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_116 =>
            -- reg_a = a2_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_117 =>
            -- reg_a = a7_X; reg_b = b1_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_118 =>
            -- reg_a = a1_X; reg_b = b7_X; reg_acc = reg_o; o8_0 = reg_o; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_119 =>
            -- reg_a = a5_X; reg_b = b4_X; reg_acc = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_120 =>
            -- reg_a = a4_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_121 =>
            -- reg_a = a6_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_122 =>
            -- reg_a = a3_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_123 =>
            -- reg_a = a7_X; reg_b = b2_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_124 =>
            -- reg_a = a2_X; reg_b = b7_X; reg_acc = reg_o; o9_0 = reg_o; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_125 =>
            -- reg_a = a5_X; reg_b = b5_X; reg_acc = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_126 =>
            -- reg_a = a6_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_127 =>
            -- reg_a = a4_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_128 =>
            -- reg_a = a7_X; reg_b = b3_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_129 =>
            -- reg_a = a3_X; reg_b = b7_X; reg_acc = reg_o; o10_0 = reg_o; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_130 =>
            -- reg_a = a6_X; reg_b = b5_X; reg_acc = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_131 =>
            -- reg_a = a5_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_132 =>
            -- reg_a = a7_X; reg_b = b4_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_133 =>
            -- reg_a = a4_X; reg_b = b7_X; reg_acc = reg_o; o11_0 = reg_o; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_134 =>
            -- reg_a = a6_X; reg_b = b6_X; reg_acc = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_135 =>
            -- reg_a = a7_X; reg_b = b5_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_136 =>
            -- reg_a = a5_X; reg_b = b7_X; reg_acc = reg_o; o12_0 = reg_o; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_137 =>
            -- reg_a = a7_X; reg_b = b6_X; reg_acc = reg_o >> 256; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_138 =>
            -- reg_a = a6_X; reg_b = b7_X; reg_acc = reg_o; o13_0 = reg_o; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_139 =>
            -- reg_a = a7_X; reg_b = b7_X; reg_acc = reg_o >> 256; o14_X = reg_o; o15_X = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_0 => 
            -- -- In case of size 1
            -- reg_a = a0_X; reg_b = a0_X; reg_acc = 0; o0_X = reg_o; o1_X = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_2 => 
            -- -- In case of sizes 2, 3, 4, 5, 6, 7, 8
            -- reg_a = a0_X; reg_b = a0_X; reg_acc = 0; o0_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_3 => 
            -- -- In case of size 2
            -- reg_a = a1_X; reg_b = a0_X; reg_acc = reg_o >> 256; o1_X = reg_o; Enable sign a; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_4 => 
            -- reg_a = a1_X; reg_b = a1_X; reg_acc = reg_o >> 256; o2_X = reg_o; o3_X = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_6 => 
            -- -- Other cases
            -- reg_a = a1_X; reg_b = a0_X; reg_acc = reg_o >> 256; o1_X = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_7 =>
            -- reg_a = a1_X; reg_b = a1_X; reg_acc = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_8 =>
            -- -- In case of size 3
            -- reg_a = a0_X; reg_b = a2_X; reg_acc = reg_o; o2_X = reg_o; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_9 =>
            -- reg_a = a2_X; reg_b = a1_X; reg_acc = reg_o >> 256; o3_X = reg_o; Enable sign a; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_10 =>
            -- reg_a = a2_X; reg_b = a2_X; reg_acc = reg_o >> 256; o4_X = reg_o; o5_X = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_12 =>
            -- -- Other cases
            -- reg_a = a0_X; reg_b = a2_X; reg_acc = reg_o; o2_X = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_13 =>
            -- reg_a = a2_X; reg_b = a1_X; reg_acc = reg_o >> 256; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_14 =>
            -- -- In case of size 4
            -- reg_a = a3_X; reg_b = a0_X; reg_acc = reg_o; o3_X = reg_o; Enable sign a; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_15 =>
            -- reg_a = a2_X; reg_b = a2_X; reg_acc = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_16 =>
            -- reg_a = a3_X; reg_b = a1_X; reg_acc = reg_o; o4_X = reg_o; Enable sign a; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_17 =>
            -- reg_a = a3_X; reg_b = a2_X; reg_acc = reg_o >> 256; o5_X = reg_o; Enable sign a; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_18 =>
            -- reg_a = a3_X; reg_b = a3_X; reg_acc = reg_o >> 256; o6_X = reg_o; o7_X = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_20 =>
            -- -- Other cases
            -- reg_a = a3_X; reg_b = a0_X; reg_acc = reg_o; o3_X = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_21 =>
            -- reg_a = a2_X; reg_b = a2_X; reg_acc = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_22 =>
            -- reg_a = a3_X; reg_b = a1_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_23 =>
            -- -- In case of size 5
            -- reg_a = a4_X; reg_b = a0_X; reg_acc = reg_o; o4_X = reg_o; Enable sign a; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_24 =>
            -- reg_a = a3_X; reg_b = a2_X; reg_acc = reg_o >> 256; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_25 =>
            -- reg_a = a4_X; reg_b = a1_X; reg_acc = reg_o; o5_X = reg_o; Enable sign a; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_26 =>
            -- reg_a = a3_X; reg_b = a3_X; reg_acc = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_27 =>
            -- reg_a = a4_X; reg_b = a2_X; reg_acc = reg_o; o6_X = reg_o; Enable sign a; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_28 =>
            -- reg_a = a4_X; reg_b = a3_X; reg_acc = reg_o >> 256; o7_X = reg_o; Enable sign a; operation : 2*a*b + acc; Increase base address o;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "111";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '1';
        when square_direct_29 =>
            -- reg_a = a4_X; reg_b = a4_X; reg_acc = reg_o >> 256; o8_X = reg_o; o9_X = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_31 =>
            -- -- Other cases
            -- reg_a = a4_X; reg_b = a0_X; reg_acc = reg_o; o4_X = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_32 =>
            -- reg_a = a3_X; reg_b = a2_X; reg_acc = reg_o >> 256; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_33 =>
            -- reg_a = a4_X; reg_b = a1_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_34 =>
            -- -- In case of size 6
            -- reg_a = a5_X; reg_b = a0_X; reg_acc = reg_o; o5_X = reg_o; Enable sign a; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_35 =>
            -- reg_a = a3_X; reg_b = a3_X; reg_acc = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_36 =>
            -- reg_a = a4_X; reg_b = a2_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_37 =>
            -- reg_a = a5_X; reg_b = a1_X; reg_acc = reg_o; o6_X = reg_o; Enable sign a; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_38 =>
            -- reg_a = a4_X; reg_b = a3_X; reg_acc = reg_o >> 256; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "111";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_39 =>
            -- reg_a = a5_X; reg_b = a2_X; reg_acc = reg_o; o7_X = reg_o; Enable sign a; operation : 2*a*b + acc; Increase base address o;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "111";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '1';
        when square_direct_40 =>
            -- reg_a = a4_X; reg_b = a4_X; reg_acc = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_41 =>
            -- reg_a = a5_X; reg_b = a3_X; reg_acc = reg_o; o8_X = reg_o; Enable sign a; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_42 =>
            -- reg_a = a5_X; reg_b = a4_X; reg_acc = reg_o >> 256; o9_X = reg_o; Enable sign a; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_43 =>
            -- reg_a = a5_X; reg_b = a5_X; reg_acc = reg_o >> 256; o10_X = reg_o; o11_X = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_45 =>
            -- -- Other cases
            -- reg_a = a5_X; reg_b = a0_X; reg_acc = reg_o; o5_X = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_46 =>
            -- reg_a = a3_X; reg_b = a3_X; reg_acc = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_47 =>
            -- reg_a = a4_X; reg_b = a2_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_48 =>
            -- reg_a = a5_X; reg_b = a1_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_49 =>
            -- -- In case of size 7
            -- reg_a = a6_X; reg_b = a0_X; reg_acc = reg_o; o6_X = reg_o; Enable sign a; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_50 =>
            -- reg_a = a4_X; reg_b = a3_X; reg_acc = reg_o >> 256; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "111";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_51 =>
            -- reg_a = a5_X; reg_b = a2_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "111";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_52 =>
            -- reg_a = a6_X; reg_b = a1_X; reg_acc = reg_o; o7_X = reg_o; Enable sign a; operation : 2*a*b + acc; Increase base address o;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "111";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '1';
        when square_direct_53 =>
            -- reg_a = a4_X; reg_b = a4_X; reg_acc = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_54 =>
            -- reg_a = a5_X; reg_b = a3_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_55 =>
            -- reg_a = a6_X; reg_b = a2_X; reg_acc = reg_o; o8_X = reg_o; Enable sign a; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_56 =>
            -- reg_a = a5_X; reg_b = a4_X; reg_acc = reg_o >> 256; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_57 =>
            -- reg_a = a6_X; reg_b = a3_X; reg_acc = reg_o; o9_X = reg_o; Enable sign a; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_58 =>
            -- reg_a = a5_X; reg_b = a5_X; reg_acc = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_59 =>
            -- reg_a = a6_X; reg_b = a4_X; reg_acc = reg_o; o10_X = reg_o; Enable sign a; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_60 =>
            -- reg_a = a6_X; reg_b = a5_X; reg_acc = reg_o >> 256; o11_X = reg_o; Enable sign a; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_61 =>
            -- reg_a = a6_X; reg_b = a6_X; reg_acc = reg_o >> 256; o12_X = reg_o; o13_X = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_63 =>
            -- -- In case of size 8
            -- reg_a = a6_X; reg_b = a0_X; reg_acc = reg_o; o6_X = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_64 =>
            -- reg_a = a4_X; reg_b = a3_X; reg_acc = reg_o >> 256; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "111";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_65 =>
            -- reg_a = a5_X; reg_b = a2_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "111";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_66 =>
            -- reg_a = a6_X; reg_b = a1_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "111";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_67 =>
            -- reg_a = a7_X; reg_b = a0_X; reg_acc = reg_o; o7_X = reg_o; Enable sign a; operation : 2*a*b + acc; Increase base address o;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "111";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '1';
        when square_direct_68 =>
            -- reg_a = a4_X; reg_b = a4_X; reg_acc = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_69 =>
            -- reg_a = a5_X; reg_b = a3_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_70 =>
            -- reg_a = a6_X; reg_b = a2_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_71 =>
            -- reg_a = a7_X; reg_b = a1_X; reg_acc = reg_o; o8_X = reg_o; Enable sign a; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_72 =>
            -- reg_a = a5_X; reg_b = a4_X; reg_acc = reg_o >> 256; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_73 =>
            -- reg_a = a6_X; reg_b = a3_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_74 =>
            -- reg_a = a7_X; reg_b = a2_X; reg_acc = reg_o; o9_X = reg_o; Enable sign a; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_75 =>
            -- reg_a = a5_X; reg_b = a5_X; reg_acc = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_76 =>
            -- reg_a = a6_X; reg_b = a4_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_77 =>
            -- reg_a = a7_X; reg_b = a3_X; reg_acc = reg_o; o10_X = reg_o; Enable sign a; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_78 =>
            -- reg_a = a6_X; reg_b = a5_X; reg_acc = reg_o >> 256; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_79 =>
            -- reg_a = a7_X; reg_b = a4_X; reg_acc = reg_o; o11_X = reg_o; Enable sign a; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_80 =>
            -- reg_a = a6_X; reg_b = a6_X; reg_acc = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_81 =>
            -- reg_a = a7_X; reg_b = a5_X; reg_acc = reg_o; o12_X = reg_o; Enable sign a; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_82 =>
            -- reg_a = a7_X; reg_b = a6_X; reg_acc = reg_o >> 256; o13_X = reg_o; Enable sign a; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_83 =>
            -- reg_a = a7_X; reg_b = a7_X; reg_acc = reg_o >> 256; o14_X = reg_o; o15_X = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
            
            
            
        when multiplication_with_reduction_0 =>
            -- -- In case of size 1
            -- reg_a = a0_X; reg_b = b0_X; reg_acc = 0; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_1 =>
            -- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o0_X = reg_y; operation : keep accumulator;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "11";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "10";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "11";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '1';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_2 =>
            -- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "01";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_3 =>
            -- reg_a = 0; reg_b = 0; reg_acc = reg_o >> 256; o0_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "11";
            next_mac_clear_reg_b <= '1';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_5 =>
            -- -- In case of sizes 2, 3, 4, 5, 6, 7, 8
            -- reg_a = a0_X; reg_b = b0_X; reg_acc = 0; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_6 =>
            -- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o0_X = reg_y; operation : keep accumulator;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "11";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "10";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "11";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '1';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_7 =>
            -- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "01";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_8 =>
            --reg_a = o0_X; reg_b = prime1; reg_acc = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_9 =>
            -- -- In case of size 2
            -- reg_a = a0_X; reg_b = b1_X; reg_acc = reg_o; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_10 =>
            -- reg_a = a1_X; reg_b = b0_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_11 =>
            -- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o1_X = reg_y; operation : keep accumulator;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "11";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "10";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "11";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '1';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_12 =>
            -- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "01";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_13 =>
            -- reg_a = a1_X; reg_b = b1_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_14 =>
            -- reg_a = o1_X; reg_b = prime1; reg_acc = reg_o; o0_X = reg_o; o1_X = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_16 =>
            -- -- Other cases
            -- reg_a = a0_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_17 =>
            -- reg_a = a1_X; reg_b = b0_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_18 =>
            -- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o1_X = reg_y; operation : keep accumulator;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "11";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "10";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "11";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '1';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_19 =>
            -- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "01";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_20 =>
            -- reg_a = o0_X; reg_b = prime2; reg_acc = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_21 =>
            -- reg_a = a1_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_22 =>
            -- reg_a = o1_X; reg_b = prime1; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_23 =>
            -- -- In case of size 3
            -- reg_a = a0_X; reg_b = b2_X; reg_acc = reg_o; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_24 =>
            -- reg_a = a2_X; reg_b = b0_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_25 =>
            -- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o2_X = reg_y; operation : keep accumulator;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "11";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "10";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "11";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '1';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_26 =>
            -- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "01";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_27 =>
            -- reg_a = a1_X; reg_b = b2_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_28 =>
            -- reg_a = o1_X; reg_b = prime2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_29 =>
            -- reg_a = a2_X; reg_b = b1_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_30 =>
            -- reg_a = o2_X; reg_b = prime1; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_31 =>
            -- reg_a = a2_X; reg_b = b2_X; reg_acc = reg_o >> 256; Enable sign a, b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_32 =>
            -- reg_a = o2_X; reg_b = prime2; reg_acc = reg_o; o1_X = reg_o; o2_X = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_34 =>
            -- -- Other cases
            -- reg_a = a0_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_35 =>
            -- reg_a = a2_X; reg_b = b0_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_36 =>
            -- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o2_X = reg_y; operation : keep accumulator;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "11";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "10";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "11";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '1';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_37 =>
            -- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "01";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_38 =>
            -- reg_a = o0_X; reg_b = prime3; reg_acc = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_39 =>
            -- reg_a = a1_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_40 =>
            -- reg_a = o1_X; reg_b = prime2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_41 =>
            -- reg_a = a2_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_42 =>
            -- reg_a = o2_X; reg_b = prime1; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_43 =>
            -- -- In case of size 4
            -- reg_a = a0_X; reg_b = b3_X; reg_acc = reg_o; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_44 =>
            -- reg_a = a3_X; reg_b = b0_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_45 =>
            -- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o3_X = reg_y; operation : keep accumulator;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "11";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "10";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "11";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '1';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_46 =>
            -- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "01";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_47 =>
            -- reg_a = a1_X; reg_b = b3_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_48 =>
            -- reg_a = o1_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_49 =>
            -- reg_a = a2_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_50 =>
            -- reg_a = o2_X; reg_b = prime2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_51 =>
            -- reg_a = a3_X; reg_b = b1_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_52 =>
            -- reg_a = o3_X; reg_b = prime1; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_53 =>
            -- reg_a = a2_X; reg_b = b3_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_54 =>
            -- reg_a = o2_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_55 =>
            -- reg_a = a3_X; reg_b = b2_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_56 =>
            -- reg_a = o3_X; reg_b = prime2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_57 =>
            -- reg_a = a3_X; reg_b = b3_X; reg_acc = reg_o >> 256; Enable sign a, b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_58 =>
            -- reg_a = o3_X; reg_b = prime3; reg_acc = reg_o; o2_X = reg_o; o3_0 = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_60 =>
            -- -- Other cases
            -- reg_a = a0_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_61 =>
            -- reg_a = a3_X; reg_b = b0_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_62 =>
            -- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o3_X = reg_y; operation : keep accumulator;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "11";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "10";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "11";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '1';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_63 =>
            -- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "01";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_64 =>
            -- reg_a = o0_X; reg_b = prime4; reg_acc = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_65 =>
            -- reg_a = a1_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_66 =>
            -- reg_a = o1_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_67 =>
            -- reg_a = a2_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_68 =>
            -- reg_a = o2_X; reg_b = prime2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_69 =>
            -- reg_a = a3_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_70 =>
            -- reg_a = o3_X; reg_b = prime1; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_71 =>
            -- -- In case of size 5
            -- reg_a = a0_X; reg_b = b4_X; reg_acc = reg_o; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_72 =>
            -- reg_a = a4_X; reg_b = b0_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_73 =>
            -- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o4_X = reg_y; operation : keep accumulator;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "11";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "10";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "11";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '1';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_74 =>
            -- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "01";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_75 =>
            -- reg_a = a1_X; reg_b = b4_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_76 =>
            -- reg_a = o1_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_77 =>
            -- reg_a = a2_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_78 =>
            -- reg_a = o2_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_79 =>
            -- reg_a = a3_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_80 =>
            -- reg_a = o3_X; reg_b = prime2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_81 =>
            -- reg_a = a4_X; reg_b = b1_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_82 =>
            -- reg_a = o4_X; reg_b = prime1; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_83 =>
            -- reg_a = a2_X; reg_b = b4_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_84 =>
            -- reg_a = o2_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_85 =>
            -- reg_a = a3_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_86 =>
            -- reg_a = o3_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_87 =>
            -- reg_a = a4_X; reg_b = b2_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_88 =>
            -- reg_a = o4_X; reg_b = prime2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_89 =>
            -- reg_a = a3_X; reg_b = b4_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_90 =>
            -- reg_a = o3_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_91 =>
            -- reg_a = a4_X; reg_b = b3_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_92 =>
            -- reg_a = o4_X; reg_b = prime3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_93 =>
            -- reg_a = a4_X; reg_b = b4_X; reg_acc = reg_o >> 256; Enable sign a, b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_94 =>
            -- reg_a = o4_X; reg_b = prime4; reg_acc = reg_o; o3_X = reg_o; o4_0 = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_96 =>
            -- -- Other cases
            -- reg_a = a0_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_97 =>
            -- reg_a = a4_X; reg_b = b0_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_98 =>
            -- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o4_X = reg_y; operation : keep accumulator;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "11";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "10";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "11";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '1';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_99 =>
            -- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "01";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_100 =>
            -- reg_a = o0_X; reg_b = prime5; reg_acc = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_101 =>
            -- reg_a = a1_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_102 =>
            -- reg_a = o1_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_103 =>
            -- reg_a = a2_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_104 =>
            -- reg_a = o2_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_105 =>
            -- reg_a = a3_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_106 =>
            -- reg_a = o3_X; reg_b = prime2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_107 =>
            -- reg_a = a4_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_108 =>
            -- reg_a = o4_X; reg_b = prime1; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_109 =>
            -- -- In case of size 6
            -- reg_a = a0_X; reg_b = b5_X; reg_acc = reg_o; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_110 =>
            -- reg_a = a5_X; reg_b = b0_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_111 =>
            -- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o5_X = reg_y; operation : keep accumulator;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "11";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "10";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "11";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '1';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_112 =>
            -- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "01";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_113 =>
            -- reg_a = a1_X; reg_b = b5_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_114 =>
            -- reg_a = o1_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_115 =>
            -- reg_a = a2_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_116 =>
            -- reg_a = o2_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_117 =>
            -- reg_a = a3_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_118 =>
            -- reg_a = o3_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_119 =>
            -- reg_a = a4_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_120 =>
            -- reg_a = o4_X; reg_b = prime2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_121 =>
            -- reg_a = a5_X; reg_b = b1_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_122 =>
            -- reg_a = o5_X; reg_b = prime1; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_123 =>
            -- reg_a = a2_X; reg_b = b5_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_124 =>
            -- reg_a = o2_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_125 =>
            -- reg_a = a3_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_126 =>
            -- reg_a = o3_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_127 =>
            -- reg_a = a4_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_128 =>
            -- reg_a = o4_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_129 =>
            -- reg_a = a5_X; reg_b = b2_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_130 =>
            -- reg_a = o5_X; reg_b = prime2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_131 =>
            -- reg_a = a3_X; reg_b = b5_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_132 =>
            -- reg_a = o3_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_133 =>
            -- reg_a = a4_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_134 =>
            -- reg_a = o4_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_135 =>
            -- reg_a = a5_X; reg_b = b3_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_136 =>
            -- reg_a = o5_X; reg_b = prime3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_137 =>
            -- reg_a = a4_X; reg_b = b5_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_138 =>
            -- reg_a = o4_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_139 =>
            -- reg_a = a5_X; reg_b = b4_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_140 =>
            -- reg_a = o5_X; reg_b = prime4; reg_acc = reg_o; o3_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_141 =>
            -- reg_a = a5_X; reg_b = b5_X; reg_acc = reg_o >> 256; Enable sign a, b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_142 =>
            -- reg_a = o5_X; reg_b = prime5; reg_acc = reg_o; o4_X = reg_o; o5_0 = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_144 =>
            -- -- Other cases
            -- reg_a = a0_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_145 =>
            -- reg_a = a5_X; reg_b = b0_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_146 =>
            -- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o5_X = reg_y; operation : keep accumulator;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "11";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "10";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "11";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '1';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_147 =>
            -- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "01";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_148 =>
            -- reg_a = o0_X; reg_b = prime6; reg_acc = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_149 =>
            -- reg_a = a1_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_150 =>
            -- reg_a = o1_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_151 =>
            -- reg_a = a2_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_152 =>
            -- reg_a = o2_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_153 =>
            -- reg_a = a3_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_154 =>
            -- reg_a = o3_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_155 =>
            -- reg_a = a4_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_156 =>
            -- reg_a = o4_X; reg_b = prime2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_157 =>
            -- reg_a = a5_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_158 =>
            -- reg_a = o5_X; reg_b = prime1; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_159 =>
            -- -- In case of size 7
            -- reg_a = a0_X; reg_b = b6_X; reg_acc = reg_o; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_160 =>
            -- reg_a = a6_X; reg_b = b0_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_161 =>
            -- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o6_X = reg_y; operation : keep accumulator;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "11";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "10";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "11";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '1';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_162 =>
            -- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "01";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_163 =>
            -- reg_a = a1_X; reg_b = b6_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_164 =>
            -- reg_a = o1_X; reg_b = prime6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_165 =>
            -- reg_a = a2_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_166 =>
            -- reg_a = o2_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_167 =>
            -- reg_a = a3_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_168 =>
            -- reg_a = o3_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_169 =>
            -- reg_a = a4_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_170 =>
            -- reg_a = o4_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_171 =>
            -- reg_a = a5_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_172 =>
            -- reg_a = o5_X; reg_b = prime2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_173 =>
            -- reg_a = a6_X; reg_b = b1_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_174 =>
            -- reg_a = o6_X; reg_b = prime1; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_175 =>
            -- reg_a = a2_X; reg_b = b6_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_176 =>
            -- reg_a = o2_X; reg_b = prime6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_177 =>
            -- reg_a = a3_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_178 =>
            -- reg_a = o3_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_179 =>
            -- reg_a = a4_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_180 =>
            -- reg_a = o4_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_181 =>
            -- reg_a = a5_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_182 =>
            -- reg_a = o5_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_183 =>
            -- reg_a = a6_X; reg_b = b2_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_184 =>
            -- reg_a = o6_X; reg_b = prime2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_185 =>
            -- reg_a = a3_X; reg_b = b6_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_186 =>
            -- reg_a = o3_X; reg_b = prime6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_187 =>
            -- reg_a = a4_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_188 =>
            -- reg_a = o4_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_189 =>
            -- reg_a = a5_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_190 =>
            -- reg_a = o5_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_191 =>
            -- reg_a = a6_X; reg_b = b3_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_192 =>
            -- reg_a = o6_X; reg_b = prime3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_193 =>
            -- reg_a = a4_X; reg_b = b6_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_194 =>
            -- reg_a = o4_X; reg_b = prime6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_195 =>
            -- reg_a = a5_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_196 =>
            -- reg_a = o5_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_197 =>
            -- reg_a = a6_X; reg_b = b4_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_198 =>
            -- reg_a = o6_X; reg_b = prime4; reg_acc = reg_o; o3_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_199 =>
            -- reg_a = a5_X; reg_b = b6_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_200 =>
            -- reg_a = o5_X; reg_b = prime6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_201 =>
            -- reg_a = a6_X; reg_b = b5_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_202 =>
            -- reg_a = o6_X; reg_b = prime5; reg_acc = reg_o; o4_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_203 =>
            -- reg_a = a6_X; reg_b = b6_X; reg_acc = reg_o >> 256; Enable sign a, b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_204 =>
            -- reg_a = o6_X; reg_b = prime6; reg_acc = reg_o; o5_X = reg_o; o6_0 = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_206 =>
            -- -- In case of size 8
            -- reg_a = a0_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_207 =>
            -- reg_a = a6_X; reg_b = b0_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_208 =>
            -- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o6_X = reg_y; operation : keep accumulator;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "11";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "10";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "11";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '1';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_209 =>
            -- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "01";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_210 =>
            -- reg_a = o0_X; reg_b = prime7; reg_acc = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_211 =>
            -- reg_a = a1_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_212 =>
            -- reg_a = o1_X; reg_b = prime6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_213 =>
            -- reg_a = a2_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_214 =>
            -- reg_a = o2_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_215 =>
            -- reg_a = a3_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_216 =>
            -- reg_a = o3_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_217 =>
            -- reg_a = a4_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_218 =>
            -- reg_a = o4_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_219 =>
            -- reg_a = a5_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_220 =>
            -- reg_a = o5_X; reg_b = prime2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_221 =>
            -- reg_a = a6_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_222 =>
            -- reg_a = o6_X; reg_b = prime1; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_223 =>
            -- reg_a = a0_X; reg_b = b7_X; reg_acc = reg_o; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_224 =>
            -- reg_a = a7_X; reg_b = b0_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_225 =>
            -- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o7_X = reg_y; operation : keep accumulator;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "11";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "111";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "10";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "11";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '1';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_226 =>
            -- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "01";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_227 =>
            -- reg_a = a1_X; reg_b = b7_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_228 =>
            -- reg_a = o1_X; reg_b = prime7; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_229 =>
            -- reg_a = a2_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_230 =>
            -- reg_a = o2_X; reg_b = prime6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_231 =>
            -- reg_a = a3_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_232 =>
            -- reg_a = o3_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_233 =>
            -- reg_a = a4_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_234 =>
            -- reg_a = o4_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_235 =>
            -- reg_a = a5_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_236 =>
            -- reg_a = o5_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_237 =>
            -- reg_a = a6_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_238 =>
            -- reg_a = o6_X; reg_b = prime2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_239 =>
            -- reg_a = a7_X; reg_b = b1_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_240 =>
            -- reg_a = o7_X; reg_b = prime1; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_241 =>
            -- reg_a = a2_X; reg_b = b7_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_242 =>
            -- reg_a = o2_X; reg_b = prime7; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_243 =>
            -- reg_a = a3_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_244 =>
            -- reg_a = o3_X; reg_b = prime6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_245 =>
            -- reg_a = a4_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_246 =>
            -- reg_a = o4_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_247 =>
            -- reg_a = a5_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_248 =>
            -- reg_a = o5_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_249 =>
            -- reg_a = a6_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_250 =>
            -- reg_a = o6_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_251 =>
            -- reg_a = a7_X; reg_b = b2_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_252 =>
            -- reg_a = o7_X; reg_b = prime2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_253 =>
            -- reg_a = a3_X; reg_b = b7_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_254 =>
            -- reg_a = o3_X; reg_b = prime7; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_255 =>
            -- reg_a = a4_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_256 =>
            -- reg_a = o4_X; reg_b = prime6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_257 =>
            -- reg_a = a5_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_258 =>
            -- reg_a = o5_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_259 =>
            -- reg_a = a6_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_260 =>
            -- reg_a = o6_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_261 =>
            -- reg_a = a7_X; reg_b = b3_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_262 =>
            -- reg_a = o7_X; reg_b = prime3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_263 =>
            -- reg_a = a4_X; reg_b = b7_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_264 =>
            -- reg_a = o4_X; reg_b = prime7; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_265 =>
            -- reg_a = a5_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_266 =>
            -- reg_a = o5_X; reg_b = prime6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_267 =>
            -- reg_a = a6_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_268 =>
            -- reg_a = o6_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_269 =>
            -- reg_a = a7_X; reg_b = b4_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_270 =>
            -- reg_a = o7_X; reg_b = prime4; reg_acc = reg_o; o3_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_271 =>
            -- reg_a = a5_X; reg_b = b7_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_272 =>
            -- reg_a = o5_X; reg_b = prime7; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_273 =>
            -- reg_a = a6_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_274 =>
            -- reg_a = o6_X; reg_b = prime6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_275 =>
            -- reg_a = a7_X; reg_b = b5_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_276 =>
            -- reg_a = o7_X; reg_b = prime5; reg_acc = reg_o; o4_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_277 =>
            -- reg_a = a6_X; reg_b = b7_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_278 =>
            -- reg_a = o6_X; reg_b = prime7; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_279 =>
            -- reg_a = a7_X; reg_b = b6_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_280 =>
            -- reg_a = o7_X; reg_b = prime6; reg_acc = reg_o; o5_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_281 =>
            -- reg_a = a7_X; reg_b = b7_X; reg_acc = reg_o >> 256; Enable sign a, b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_282 =>
            -- reg_a = o7_X; reg_b = prime7; reg_acc = reg_o; o6_X = reg_o; o7_0 = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_0 =>
            -- -- In case of size 1
            -- reg_a = a0_X; reg_b = b0_X; reg_acc = 0; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_1 =>
            -- reg_a = 0; reg_b = 0; reg_acc = reg_o >> 256; o0_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "11";
            next_mac_clear_reg_b <= '1';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_3 =>
            -- -- In case of sizes 2, 3, 4, 5, 6, 7, 8
            -- reg_a = a0_X; reg_b = b0_X; reg_acc = 0; o0_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_4 =>
            -- -- In case of size 2
            -- reg_a = a0_X; reg_b = b1_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_5 =>
            -- reg_a = o0_X; reg_b = primeSP1; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_6 =>
            -- reg_a = a1_X; reg_b = b0_X; reg_acc = reg_o; o1_X = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_7 =>
            -- reg_a = a1_X; reg_b = b1_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_8 =>
            -- reg_a = o1_X; reg_b = primeSP1; reg_acc = reg_o; o0_X = reg_o; o1_X = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_10 =>
            -- -- In case of sizes 3, 4, 5, 6, 7, 8
            -- reg_a = a0_X; reg_b = b1_X; reg_acc = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_11 =>
            -- reg_a = o0_X; reg_b = primeSP1; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_12 =>
            -- reg_a = a1_X; reg_b = b0_X; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_13 =>
            -- reg_a = o0_X; reg_b = primeSP2; reg_acc = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_14 =>
            -- reg_a = a1_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_15 =>
            -- reg_a = o1_X; reg_b = primeSP1; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_16 =>
            -- -- In case of size 3
            -- reg_a = a0_X; reg_b = b2_X; reg_acc = reg_o; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_17 =>
            -- reg_a = a2_X; reg_b = b0_X; reg_acc = reg_o; o2_X = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_18 =>
            -- reg_a = a1_X; reg_b = b2_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_19 =>
            -- reg_a = o1_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_20 =>
            -- reg_a = a2_X; reg_b = b1_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_21 =>
            -- reg_a = o2_X; reg_b = primeSP1; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_22 =>
            -- reg_a = a2_X; reg_b = b2_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_23 =>
            -- reg_a = o2_X; reg_b = primeSP2; reg_acc = reg_o; o1_X = reg_o; o2_X = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_25 =>
            -- -- In case of sizes 4, 5, 6, 7, 8
            -- reg_a = a0_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_26 =>
            -- reg_a = a2_X; reg_b = b0_X; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_27 =>
            -- reg_a = o0_X; reg_b = primeSP3; reg_acc = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_28 =>
            -- reg_a = a1_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_29 =>
            -- reg_a = o1_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_30 =>
            -- reg_a = a2_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_31 =>
            -- reg_a = o2_X; reg_b = primeSP1; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_32 =>
            -- -- In case of size 4
            -- reg_a = a0_X; reg_b = b3_X; reg_acc = reg_o; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_33 =>
            -- reg_a = a3_X; reg_b = b0_X; reg_acc = reg_o; o3_X = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_34 =>
            -- reg_a = a1_X; reg_b = b3_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_35 =>
            -- reg_a = o1_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_36 =>
            -- reg_a = a2_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_37 =>
            -- reg_a = o2_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_38 =>
            -- reg_a = a3_X; reg_b = b1_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_39 =>
            -- reg_a = o3_X; reg_b = primeSP1; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_40 =>
            -- reg_a = a2_X; reg_b = b3_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_41 =>
            -- reg_a = o2_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_42 =>
            -- reg_a = a3_X; reg_b = b2_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_43 =>
            -- reg_a = o3_X; reg_b = primeSP2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_44 =>
            -- reg_a = a3_X; reg_b = b3_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_45 =>
            -- reg_a = o3_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; o3_X = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_47 =>
            -- -- In case of sizes 5, 6, 7, 8
            -- reg_a = a0_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_48 =>
            -- reg_a = a3_X; reg_b = b0_X; reg_acc = reg_o; o3_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_49 =>
            -- reg_a = o0_X; reg_b = primeSP4; reg_acc = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_50 =>
            -- reg_a = a1_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_51 =>
            -- reg_a = o1_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_52 =>
            -- reg_a = a2_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_53 =>
            -- reg_a = o2_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_54 =>
            -- reg_a = a3_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_55 =>
            -- reg_a = o3_X; reg_b = primeSP1; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_56 =>
            -- -- In case of size 5
            -- reg_a = a0_X; reg_b = b4_X; reg_acc = reg_o; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_57 =>
            -- reg_a = a4_X; reg_b = b0_X; reg_acc = reg_o; o4_X = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_58 =>
            -- reg_a = a1_X; reg_b = b4_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_59 =>
            -- reg_a = o1_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_60 =>
            -- reg_a = a2_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_61 =>
            -- reg_a = o2_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_62 =>
            -- reg_a = a3_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_63 =>
            -- reg_a = o3_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_64 =>
            -- reg_a = a4_X; reg_b = b1_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_65 =>
            -- reg_a = o4_X; reg_b = primeSP1; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_66 =>
            -- reg_a = a2_X; reg_b = b4_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_67 =>
            -- reg_a = o2_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_68 =>
            -- reg_a = a3_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_69 =>
            -- reg_a = o3_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_70 =>
            -- reg_a = a4_X; reg_b = b2_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_71 =>
            -- reg_a = o4_X; reg_b = primeSP2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_72 =>
            -- reg_a = a3_X; reg_b = b4_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_73 =>
            -- reg_a = o3_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_74 =>
            -- reg_a = a4_X; reg_b = b3_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_75 =>
            -- reg_a = o4_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_76 =>
            -- reg_a = a4_X; reg_b = b4_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_77 =>
            -- reg_a = o4_X; reg_b = primeSP4; reg_acc = reg_o; o3_X = reg_o; o4_X = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_79 =>
            -- -- In case of sizes 6, 7, 8
            -- reg_a = a0_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_80 =>
            -- reg_a = a4_X; reg_b = b0_X; reg_acc = reg_o; o4_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_81 =>
            -- reg_a = o0_X; reg_b = primeSP5; reg_acc = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_82 =>
            -- reg_a = a1_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_83 =>
            -- reg_a = o1_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_84 =>
            -- reg_a = a2_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_85 =>
            -- reg_a = o2_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_86 =>
            -- reg_a = a3_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_87 =>
            -- reg_a = o3_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_88 =>
            -- reg_a = a4_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_89 =>
            -- reg_a = o4_X; reg_b = primeSP1; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_90 =>
            -- -- In case of size 6
            -- reg_a = a0_X; reg_b = b5_X; reg_acc = reg_o; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_91 =>
            -- reg_a = a5_X; reg_b = b0_X; reg_acc = reg_o; o5_X = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_92 =>
            -- reg_a = a1_X; reg_b = b5_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_93 =>
            -- reg_a = o1_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_94 =>
            -- reg_a = a2_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_95 =>
            -- reg_a = o2_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_96 =>
            -- reg_a = a3_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_97 =>
            -- reg_a = o3_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_98 =>
            -- reg_a = a4_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_99 =>
            -- reg_a = o4_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_100 =>
            -- reg_a = a5_X; reg_b = b1_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_101 =>
            -- reg_a = o5_X; reg_b = primeSP1; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_102 =>
            -- reg_a = a2_X; reg_b = b5_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_103 =>
            -- reg_a = o2_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_104 =>
            -- reg_a = a3_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_105 =>
            -- reg_a = o3_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_106 =>
            -- reg_a = a4_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_107 =>
            -- reg_a = o4_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_108 =>
            -- reg_a = a5_X; reg_b = b2_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_109 =>
            -- reg_a = o5_X; reg_b = primeSP2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_110 =>
            -- reg_a = a3_X; reg_b = b5_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_111 =>
            -- reg_a = o3_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_112 =>
            -- reg_a = a4_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_113 =>
            -- reg_a = o4_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_114 =>
            -- reg_a = a5_X; reg_b = b3_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_115 =>
            -- reg_a = o5_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_116 =>
            -- reg_a = a4_X; reg_b = b5_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_117 =>
            -- reg_a = o4_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_118 =>
            -- reg_a = a5_X; reg_b = b4_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_119 =>
            -- reg_a = o5_X; reg_b = primeSP4; reg_acc = reg_o; o3_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_120 =>
            -- reg_a = a5_X; reg_b = b5_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_121 =>
            -- reg_a = o5_X; reg_b = primeSP5; reg_acc = reg_o; o4_X = reg_o; o5_X = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_123 =>
            -- -- In case of sizes 7, 8
            -- reg_a = a0_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_124 =>
            -- reg_a = a5_X; reg_b = b0_X; reg_acc = reg_o; o5_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_125 =>
            -- reg_a = o0_X; reg_b = primeSP6; reg_acc = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_126 =>
            -- reg_a = a1_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_127 =>
            -- reg_a = o1_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_128 =>
            -- reg_a = a2_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_129 =>
            -- reg_a = o2_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_130 =>
            -- reg_a = a3_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_131 =>
            -- reg_a = o3_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_132 =>
            -- reg_a = a4_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_133 =>
            -- reg_a = o4_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_134 =>
            -- reg_a = a5_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_135 =>
            -- reg_a = o5_X; reg_b = primeSP1; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_136 =>
            -- -- In case of size 7
            -- reg_a = a0_X; reg_b = b6_X; reg_acc = reg_o; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_137 =>
            -- reg_a = a6_X; reg_b = b0_X; reg_acc = reg_o; o6_X = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_138 =>
            -- reg_a = a1_X; reg_b = b6_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_139 =>
            -- reg_a = o1_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_140 =>
            -- reg_a = a2_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_141 =>
            -- reg_a = o2_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_142 =>
            -- reg_a = a3_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_143 =>
            -- reg_a = o3_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_144 =>
            -- reg_a = a4_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_145 =>
            -- reg_a = o4_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_146 =>
            -- reg_a = a5_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_147 =>
            -- reg_a = o5_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_148 =>
            -- reg_a = a6_X; reg_b = b1_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_149 =>
            -- reg_a = o6_X; reg_b = primeSP1; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_150 =>
            -- reg_a = a2_X; reg_b = b6_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_151 =>
            -- reg_a = o2_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_152 =>
            -- reg_a = a3_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_153 =>
            -- reg_a = o3_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_154 =>
            -- reg_a = a4_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_155 =>
            -- reg_a = o4_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_156 =>
            -- reg_a = a5_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_157 =>
            -- reg_a = o5_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_158 =>
            -- reg_a = a6_X; reg_b = b2_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_159 =>
            -- reg_a = o6_X; reg_b = primeSP2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_160 =>
            -- reg_a = a3_X; reg_b = b6_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_161 =>
            -- reg_a = o3_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_162 =>
            -- reg_a = a4_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_163 =>
            -- reg_a = o4_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_164 =>
            -- reg_a = a5_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_165 =>
            -- reg_a = o5_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_166 =>
            -- reg_a = a6_X; reg_b = b3_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_167 =>
            -- reg_a = o6_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_168 =>
            -- reg_a = a4_X; reg_b = b6_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_169 =>
            -- reg_a = o4_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_170 =>
            -- reg_a = a5_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_171 =>
            -- reg_a = o5_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_172 =>
            -- reg_a = a6_X; reg_b = b4_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_173 =>
            -- reg_a = o6_X; reg_b = primeSP4; reg_acc = reg_o; o3_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_174 =>
            -- reg_a = a5_X; reg_b = b6_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_175 =>
            -- reg_a = o5_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_176 =>
            -- reg_a = a6_X; reg_b = b5_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_177 =>
            -- reg_a = o6_X; reg_b = primeSP5; reg_acc = reg_o; o4_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_178 =>
            -- reg_a = a6_X; reg_b = b6_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_179 =>
            -- reg_a = o6_X; reg_b = primeSP6; reg_acc = reg_o; o5_X = reg_o; o6_X = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_181 =>
            -- -- In case of size 8
            -- reg_a = a0_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_182 =>
            -- reg_a = a6_X; reg_b = b0_X; reg_acc = reg_o; o6_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_183 =>
            -- reg_a = o0_X; reg_b = primeSP7; reg_acc = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_184 =>
            -- reg_a = a1_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_185 =>
            -- reg_a = o1_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_186 =>
            -- reg_a = a2_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_187 =>
            -- reg_a = o2_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_188 =>
            -- reg_a = a3_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_189 =>
            -- reg_a = o3_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_190 =>
            -- reg_a = a4_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_191 =>
            -- reg_a = o4_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_192 =>
            -- reg_a = a5_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_193 =>
            -- reg_a = o5_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_194 =>
            -- reg_a = a6_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_195 =>
            -- reg_a = o6_X; reg_b = primeSP1; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_196 =>
            -- reg_a = a0_X; reg_b = b7_X; reg_acc = reg_o; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_197 =>
            -- reg_a = a7_X; reg_b = b0_X; reg_acc = reg_o; o7_X = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "111";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_198 =>
            -- reg_a = a1_X; reg_b = b7_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_199 =>
            -- reg_a = o1_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_200 =>
            -- reg_a = a2_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_201 =>
            -- reg_a = o2_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_202 =>
            -- reg_a = a3_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_203 =>
            -- reg_a = o3_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_204 =>
            -- reg_a = a4_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_205 =>
            -- reg_a = o4_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_206 =>
            -- reg_a = a5_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_207 =>
            -- reg_a = o5_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_208 =>
            -- reg_a = a6_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_209 =>
            -- reg_a = o6_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_210 =>
            -- reg_a = a7_X; reg_b = b1_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_211 =>
            -- reg_a = o7_X; reg_b = primeSP1; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_212 =>
            -- reg_a = a2_X; reg_b = b7_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_213 =>
            -- reg_a = o2_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_214 =>
            -- reg_a = a3_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_215 =>
            -- reg_a = o3_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_216 =>
            -- reg_a = a4_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_217 =>
            -- reg_a = o4_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_218 =>
            -- reg_a = a5_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_219 =>
            -- reg_a = o5_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_220 =>
            -- reg_a = a6_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_221 =>
            -- reg_a = o6_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_222 =>
            -- reg_a = a7_X; reg_b = b2_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_223 =>
            -- reg_a = o7_X; reg_b = primeSP2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_224 =>
            -- reg_a = a3_X; reg_b = b7_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_225 =>
            -- reg_a = o3_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_226 =>
            -- reg_a = a4_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_227 =>
            -- reg_a = o4_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_228 =>
            -- reg_a = a5_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_229 =>
            -- reg_a = o5_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_230 =>
            -- reg_a = a6_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_231 =>
            -- reg_a = o6_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_232 =>
            -- reg_a = a7_X; reg_b = b3_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_233 =>
            -- reg_a = o7_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_234 =>
            -- reg_a = a4_X; reg_b = b7_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_235 =>
            -- reg_a = o4_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_236 =>
            -- reg_a = a5_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_237 =>
            -- reg_a = o5_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_238 =>
            -- reg_a = a6_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_239 =>
            -- reg_a = o6_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_240 =>
            -- reg_a = a7_X; reg_b = b4_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_241 =>
            -- reg_a = o7_X; reg_b = primeSP4; reg_acc = reg_o; o3_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_242 =>
            -- reg_a = a5_X; reg_b = b7_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_243 =>
            -- reg_a = o5_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_244 =>
            -- reg_a = a6_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_245 =>
            -- reg_a = o6_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_246 =>
            -- reg_a = a7_X; reg_b = b5_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_247 =>
            -- reg_a = o7_X; reg_b = primeSP5; reg_acc = reg_o; o4_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_248 =>
            -- reg_a = a6_X; reg_b = b7_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_249 =>
            -- reg_a = o6_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_250 =>
            -- reg_a = a7_X; reg_b = b6_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_251 =>
            -- reg_a = o7_X; reg_b = primeSP6; reg_acc = reg_o; o5_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_252 =>
            -- reg_a = a7_X; reg_b = b7_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_253 =>
            -- reg_a = o7_X; reg_b = primeSP7; reg_acc = reg_o; o6_X = reg_o; o7_X = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_0 =>
            -- With 2 zeroes in prime sharp
            -- -- In case of sizes 2, 3, 4, 5, 6, 7, 8
            -- reg_a = a0_X; reg_b = b0_X; reg_acc = 0; o0_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_1 =>
            -- -- In case of size 2
            -- reg_a = a0_X; reg_b = b1_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_2 =>
            -- reg_a = a1_X; reg_b = b0_X; reg_acc = reg_o; o1_X = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_3 =>
            -- reg_a = a1_X; reg_b = b1_X; reg_acc = reg_o >> 256; o0_X = reg_o; o1_X = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_5 =>
            -- -- In case of sizes 3, 4, 5, 6, 7, 8
            -- reg_a = a0_X; reg_b = b1_X; reg_acc = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_6 =>
            -- reg_a = a1_X; reg_b = b0_X; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_7 =>
            -- reg_a = o0_X; reg_b = primeSP2; reg_acc = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_8 =>
            -- reg_a = a1_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_9 =>
            -- -- In case of size 3
            -- reg_a = a0_X; reg_b = b2_X; reg_acc = reg_o; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_10 =>
            -- reg_a = a2_X; reg_b = b0_X; reg_acc = reg_o; o2_X = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_11 =>
            -- reg_a = a1_X; reg_b = b2_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_12 =>
            -- reg_a = o1_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_13 =>
            -- reg_a = a2_X; reg_b = b1_X; reg_acc = reg_o; Enable sign a; o0_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_14 =>
            -- reg_a = a2_X; reg_b = b2_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_15 =>
            -- reg_a = o2_X; reg_b = primeSP2; reg_acc = reg_o; o1_X = reg_o; o2_X = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_17 =>
            -- -- In case of sizes 4, 5, 6, 7, 8
            -- reg_a = a0_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_18 =>
            -- reg_a = a2_X; reg_b = b0_X; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_19 =>
            -- reg_a = o0_X; reg_b = primeSP3; reg_acc = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_20 =>
            -- reg_a = a1_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_21 =>
            -- reg_a = o1_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_22 =>
            -- reg_a = a2_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_23 =>
            -- -- In case of size 4
            -- reg_a = a0_X; reg_b = b3_X; reg_acc = reg_o; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_24 =>
            -- reg_a = a3_X; reg_b = b0_X; reg_acc = reg_o; o3_X = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_25 =>
            -- reg_a = a1_X; reg_b = b3_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_26 =>
            -- reg_a = o1_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_27 =>
            -- reg_a = a2_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_28 =>
            -- reg_a = o2_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_29 =>
            -- reg_a = a3_X; reg_b = b1_X; reg_acc = reg_o; Enable sign a; o0_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_30 =>
            -- reg_a = a2_X; reg_b = b3_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_31 =>
            -- reg_a = o2_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_32 =>
            -- reg_a = a3_X; reg_b = b2_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_33 =>
            -- reg_a = o3_X; reg_b = primeSP2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_34 =>
            -- reg_a = a3_X; reg_b = b3_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_35 =>
            -- reg_a = o3_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; o3_X = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_37 =>
            -- -- In case of sizes 5, 6, 7, 8
            -- reg_a = a0_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_38 =>
            -- reg_a = a3_X; reg_b = b0_X; reg_acc = reg_o; o3_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_39 =>
            -- reg_a = o0_X; reg_b = primeSP4; reg_acc = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_40 =>
            -- reg_a = a1_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_41 =>
            -- reg_a = o1_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_42 =>
            -- reg_a = a2_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_43 =>
            -- reg_a = o2_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_44 =>
            -- reg_a = a3_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_45 =>
            -- In case of size 5
            -- reg_a = a0_X; reg_b = b4_X; reg_acc = reg_o; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_46 =>
            -- reg_a = a4_X; reg_b = b0_X; reg_acc = reg_o; o4_X = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_47 =>
            -- reg_a = a1_X; reg_b = b4_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_48 =>
            -- reg_a = o1_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_49 =>
            -- reg_a = a2_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_50 =>
            -- reg_a = o2_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_51 =>
            -- reg_a = a3_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_52 =>
            -- reg_a = o3_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_53 =>
            -- reg_a = a4_X; reg_b = b1_X; reg_acc = reg_o; o0_X = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_54 =>
            -- reg_a = a2_X; reg_b = b4_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_55 =>
            -- reg_a = o2_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_56 =>
            -- reg_a = a3_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_57 =>
            -- reg_a = o3_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_58 =>
            -- reg_a = a4_X; reg_b = b2_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_59 =>
            -- reg_a = o4_X; reg_b = primeSP2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_60 =>
            -- reg_a = a3_X; reg_b = b4_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_61 =>
            -- reg_a = o3_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_62 =>
            -- reg_a = a4_X; reg_b = b3_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_63 =>
            -- reg_a = o4_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_64 =>
            -- reg_a = a4_X; reg_b = b4_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_65 =>
            -- reg_a = o4_X; reg_b = primeSP4; reg_acc = reg_o; o3_X = reg_o; o4_X = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_67 =>
            -- -- In case of sizes 6, 7, 8
            -- reg_a = a0_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_68 =>
            -- reg_a = a4_X; reg_b = b0_X; reg_acc = reg_o; o4_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_69 =>
            -- reg_a = o0_X; reg_b = primeSP5; reg_acc = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_70 =>
            -- reg_a = a1_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_71 =>
            -- reg_a = o1_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_72 =>
            -- reg_a = a2_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_73 =>
            -- reg_a = o2_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_74 =>
            -- reg_a = a3_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_75 =>
            -- reg_a = o3_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_76 =>
            -- reg_a = a4_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_77 =>
            -- In case of size 6
            -- reg_a = a0_X; reg_b = b5_X; reg_acc = reg_o; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_78 =>
            -- reg_a = a5_X; reg_b = b0_X; reg_acc = reg_o; o5_X = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_79 =>
            -- reg_a = a1_X; reg_b = b5_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_80 =>
            -- reg_a = o1_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_81 =>
            -- reg_a = a2_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_82 =>
            -- reg_a = o2_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_83 =>
            -- reg_a = a3_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_84 =>
            -- reg_a = o3_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_85 =>
            -- reg_a = a4_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_86 =>
            -- reg_a = o4_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_87 =>
            -- reg_a = a5_X; reg_b = b1_X; reg_acc = reg_o; o0_X = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_88 =>
            -- reg_a = a2_X; reg_b = b5_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_89 =>
            -- reg_a = o2_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_90 =>
            -- reg_a = a3_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_91 =>
            -- reg_a = o3_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_92 =>
            -- reg_a = a4_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_93 =>
            -- reg_a = o4_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_94 =>
            -- reg_a = a5_X; reg_b = b2_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_95 =>
            -- reg_a = o5_X; reg_b = primeSP2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_96 =>
            -- reg_a = a3_X; reg_b = b5_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_97 =>
            -- reg_a = o3_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_98 =>
            -- reg_a = a4_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_99 =>
            -- reg_a = o4_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_100 =>
            -- reg_a = a5_X; reg_b = b3_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_101 =>
            -- reg_a = o5_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_102 =>
            -- reg_a = a4_X; reg_b = b5_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_103 =>
            -- reg_a = o4_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_104 =>
            -- reg_a = a5_X; reg_b = b4_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_105 =>
            -- reg_a = o5_X; reg_b = primeSP4; reg_acc = reg_o; o3_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_106 =>
            -- reg_a = a5_X; reg_b = b5_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_107 =>
            -- reg_a = o5_X; reg_b = primeSP5; reg_acc = reg_o; o4_X = reg_o; o5_X = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_109 =>
            -- -- In case of sizes 7, 8
            -- reg_a = a0_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_110 =>
            -- reg_a = a5_X; reg_b = b0_X; reg_acc = reg_o; o5_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_111 =>
            -- reg_a = o0_X; reg_b = primeSP6; reg_acc = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_112 =>
            -- reg_a = a1_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_113 =>
            -- reg_a = o1_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_114 =>
            -- reg_a = a2_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_115 =>
            -- reg_a = o2_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_116 =>
            -- reg_a = a3_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_117 =>
            -- reg_a = o3_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_118 =>
            -- reg_a = a4_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_119 =>
            -- reg_a = o4_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_120 =>
            -- reg_a = a5_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_121 =>
            -- -- In case of size 7
            -- reg_a = a0_X; reg_b = b6_X; reg_acc = reg_o; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_122 =>
            -- reg_a = a6_X; reg_b = b0_X; reg_acc = reg_o; o6_X = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_123 =>
            -- reg_a = a1_X; reg_b = b6_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_124 =>
            -- reg_a = o1_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_125 =>
            -- reg_a = a2_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_126 =>
            -- reg_a = o2_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_127 =>
            -- reg_a = a3_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_128 =>
            -- reg_a = o3_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_129 =>
            -- reg_a = a4_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_130 =>
            -- reg_a = o4_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_131 =>
            -- reg_a = a5_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_132 =>
            -- reg_a = o5_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_133 =>
            -- reg_a = a6_X; reg_b = b1_X; reg_acc = reg_o; Enable sign a; o0_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_134 =>
            -- reg_a = a2_X; reg_b = b6_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_135 =>
            -- reg_a = o2_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_136 =>
            -- reg_a = a3_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_137 =>
            -- reg_a = o3_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_138 =>
            -- reg_a = a4_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_139 =>
            -- reg_a = o4_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_140 =>
            -- reg_a = a5_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_141 =>
            -- reg_a = o5_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_142 =>
            -- reg_a = a6_X; reg_b = b2_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_143 =>
            -- reg_a = o6_X; reg_b = primeSP2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_144 =>
            -- reg_a = a3_X; reg_b = b6_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_145 =>
            -- reg_a = o3_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_146 =>
            -- reg_a = a4_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_147 =>
            -- reg_a = o4_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_148 =>
            -- reg_a = a5_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_149 =>
            -- reg_a = o5_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_150 =>
            -- reg_a = a6_X; reg_b = b3_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_151 =>
            -- reg_a = o6_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_152 =>
            -- reg_a = a4_X; reg_b = b6_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_153 =>
            -- reg_a = o4_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_154 =>
            -- reg_a = a5_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_155 =>
            -- reg_a = o5_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_156 =>
            -- reg_a = a6_X; reg_b = b4_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_157 =>
            -- reg_a = o6_X; reg_b = primeSP4; reg_acc = reg_o; o3_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_158 =>
            -- reg_a = a5_X; reg_b = b6_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_159 =>
            -- reg_a = o5_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_160 =>
            -- reg_a = a6_X; reg_b = b5_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_161 =>
            -- reg_a = o6_X; reg_b = primeSP5; reg_acc = reg_o; o4_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_162 =>
            -- reg_a = a6_X; reg_b = b6_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_163 =>
            -- reg_a = o6_X; reg_b = primeSP6; reg_acc = reg_o; o5_X = reg_o; o6_X = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_165 =>
            -- -- In case of size 8
            -- reg_a = a0_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_166 =>
            -- reg_a = a6_X; reg_b = b0_X; reg_acc = reg_o; o6_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_167 =>
            -- reg_a = o0_X; reg_b = primeSP7; reg_acc = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_168 =>
            -- reg_a = a1_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_169 =>
            -- reg_a = o1_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_170 =>
            -- reg_a = a2_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_171 =>
            -- reg_a = o2_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_172 =>
            -- reg_a = a3_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_173 =>
            -- reg_a = o3_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_174 =>
            -- reg_a = a4_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_175 =>
            -- reg_a = o4_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_176 =>
            -- reg_a = a5_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_177 =>
            -- reg_a = o5_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_178 =>
            -- reg_a = a6_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_179 =>
            -- reg_a = a0_X; reg_b = b7_X; reg_acc = reg_o; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_180 =>
            -- reg_a = a7_X; reg_b = b0_X; reg_acc = reg_o; o7_X = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "111";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_181 =>
            -- reg_a = a1_X; reg_b = b7_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_182 =>
            -- reg_a = o1_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_183 =>
            -- reg_a = a2_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_184 =>
            -- reg_a = o2_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_185 =>
            -- reg_a = a3_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_186 =>
            -- reg_a = o3_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_187 =>
            -- reg_a = a4_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_188 =>
            -- reg_a = o4_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_189 =>
            -- reg_a = a5_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_190 =>
            -- reg_a = o5_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_191 =>
            -- reg_a = a6_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_192 =>
            -- reg_a = o6_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_193 =>
            -- reg_a = a7_X; reg_b = b1_X; reg_acc = reg_o; Enable sign a; o0_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_194 =>
            -- reg_a = a2_X; reg_b = b7_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_195 =>
            -- reg_a = o2_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_196 =>
            -- reg_a = a3_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_197 =>
            -- reg_a = o3_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_198 =>
            -- reg_a = a4_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_199 =>
            -- reg_a = o4_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_200 =>
            -- reg_a = a5_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_201 =>
            -- reg_a = o5_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_202 =>
            -- reg_a = a6_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_203 =>
            -- reg_a = o6_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_204 =>
            -- reg_a = a7_X; reg_b = b2_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_205 =>
            -- reg_a = o7_X; reg_b = primeSP2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_206 =>
            -- reg_a = a3_X; reg_b = b7_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_207 =>
            -- reg_a = o3_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_208 =>
            -- reg_a = a4_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_209 =>
            -- reg_a = o4_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_210 =>
            -- reg_a = a5_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_211 =>
            -- reg_a = o5_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_212 =>
            -- reg_a = a6_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_213 =>
            -- reg_a = o6_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_214 =>
            -- reg_a = a7_X; reg_b = b3_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_215 =>
            -- reg_a = o7_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_216 =>
            -- reg_a = a4_X; reg_b = b7_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_217 =>
            -- reg_a = o4_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_218 =>
            -- reg_a = a5_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_219 =>
            -- reg_a = o5_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_220 =>
            -- reg_a = a6_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_221 =>
            -- reg_a = o6_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_222 =>
            -- reg_a = a7_X; reg_b = b4_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_223 =>
            -- reg_a = o7_X; reg_b = primeSP4; reg_acc = reg_o; o3_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_224 =>
            -- reg_a = a5_X; reg_b = b7_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_225 =>
            -- reg_a = o5_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_226 =>
            -- reg_a = a6_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_227 =>
            -- reg_a = o6_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_228 =>
            -- reg_a = a7_X; reg_b = b5_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_229 =>
            -- reg_a = o7_X; reg_b = primeSP5; reg_acc = reg_o; o4_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_230 =>
            -- reg_a = a6_X; reg_b = b7_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_231 =>
            -- reg_a = o6_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_232 =>
            -- reg_a = a7_X; reg_b = b6_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_233 =>
            -- reg_a = o7_X; reg_b = primeSP6; reg_acc = reg_o; o5_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_234 =>
            -- reg_a = a7_X; reg_b = b7_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_235 =>
            -- reg_a = o7_X; reg_b = primeSP7; reg_acc = reg_o; o6_X = reg_o; o7_X = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_0 =>
            -- -- In case of sizes 3, 4, 5, 6, 7, 8
            -- reg_a = a0_X; reg_b = b0_X; reg_acc = 0; o0_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_1 =>
            -- reg_a = a0_X; reg_b = b1_X; reg_acc = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_2 =>
            -- reg_a = a1_X; reg_b = b0_X; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_3 =>
            -- reg_a = a1_X; reg_b = b1_X; reg_acc = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_4 =>
            -- -- In case of size 3
            -- reg_a = a0_X; reg_b = b2_X; reg_acc = reg_o; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_5 =>
            -- reg_a = a2_X; reg_b = b0_X; reg_acc = reg_o; o2_X = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_6 =>
            -- reg_a = a1_X; reg_b = b2_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_7 =>
            -- reg_a = a2_X; reg_b = b1_X; reg_acc = reg_o; Enable sign a; o0_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_8 =>
            -- reg_a = a2_X; reg_b = b2_X; reg_acc = reg_o >> 256; Enable sign a,b; o1_X = reg_o; o2_X = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_10 =>
            -- -- In case of sizes 4, 5, 6, 7, 8
            -- reg_a = a0_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_11 =>
            -- reg_a = a2_X; reg_b = b0_X; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_12 =>
            -- reg_a = o0_X; reg_b = primeSP3; reg_acc = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_13 =>
            -- reg_a = a1_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_14 =>
            -- reg_a = a2_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_15 =>
            -- -- In case of size 4
            -- reg_a = a0_X; reg_b = b3_X; reg_acc = reg_o; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_16 =>
            -- reg_a = a3_X; reg_b = b0_X; reg_acc = reg_o; o3_X = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_17 =>
            -- reg_a = a1_X; reg_b = b3_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_18 =>
            -- reg_a = o1_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_19 =>
            -- reg_a = a2_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_20 =>
            -- reg_a = a3_X; reg_b = b1_X; reg_acc = reg_o; Enable sign a; o0_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_21 =>
            -- reg_a = a2_X; reg_b = b3_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_22 =>
            -- reg_a = o2_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_23 =>
            -- reg_a = a3_X; reg_b = b2_X; reg_acc = reg_o; Enable sign a; o1_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_24 =>
            -- reg_a = a3_X; reg_b = b3_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_25 =>
            -- reg_a = o3_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; o3_X = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_27 =>
            -- -- In case of sizes 5, 6, 7, 8
            -- reg_a = a0_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_28 =>
            -- reg_a = a3_X; reg_b = b0_X; reg_acc = reg_o; o3_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_29 =>
            -- reg_a = o0_X; reg_b = primeSP4; reg_acc = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_30 =>
            -- reg_a = a1_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_31 =>
            -- reg_a = o1_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_32 =>
            -- reg_a = a2_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_33 =>
            -- reg_a = a3_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_34 =>
            -- In case of size 5
            -- reg_a = a0_X; reg_b = b4_X; reg_acc = reg_o; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_35 =>
            -- reg_a = a4_X; reg_b = b0_X; reg_acc = reg_o; o4_X = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_36 =>
            -- reg_a = a1_X; reg_b = b4_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_37 =>
            -- reg_a = o1_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_38 =>
            -- reg_a = a2_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_39 =>
            -- reg_a = o2_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_40 =>
            -- reg_a = a3_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_41 =>
            -- reg_a = a4_X; reg_b = b1_X; reg_acc = reg_o; o0_X = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_42 =>
            -- reg_a = a2_X; reg_b = b4_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_43 =>
            -- reg_a = o2_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_44 =>
            -- reg_a = a3_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_45 =>
            -- reg_a = o3_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_46 =>
            -- reg_a = a4_X; reg_b = b2_X; reg_acc = reg_o; Enable sign a; o1_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_47 =>
            -- reg_a = a3_X; reg_b = b4_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_48 =>
            -- reg_a = o3_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_49 =>
            -- reg_a = a4_X; reg_b = b3_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_50 =>
            -- reg_a = o4_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_51 =>
            -- reg_a = a4_X; reg_b = b4_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_52 =>
            -- reg_a = o4_X; reg_b = primeSP4; reg_acc = reg_o; o3_X = reg_o; o4_X = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_54 =>
            -- -- In case of sizes 6, 7, 8
            -- reg_a = a0_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_55 =>
            -- reg_a = a4_X; reg_b = b0_X; reg_acc = reg_o; o4_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_56 =>
            -- reg_a = o0_X; reg_b = primeSP5; reg_acc = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_57 =>
            -- reg_a = a1_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_58 =>
            -- reg_a = o1_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_59 =>
            -- reg_a = a2_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_60 =>
            -- reg_a = o2_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_61 =>
            -- reg_a = a3_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_62 =>
            -- reg_a = a4_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_63 =>
            -- In case of size 6
            -- reg_a = a0_X; reg_b = b5_X; reg_acc = reg_o; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_64 =>
            -- reg_a = a5_X; reg_b = b0_X; reg_acc = reg_o; o5_X = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_65 =>
            -- reg_a = a1_X; reg_b = b5_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_66 =>
            -- reg_a = o1_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_67 =>
            -- reg_a = a2_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_68 =>
            -- reg_a = o2_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_69 =>
            -- reg_a = a3_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_70 =>
            -- reg_a = o3_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_71 =>
            -- reg_a = a4_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_72 =>
            -- reg_a = a5_X; reg_b = b1_X; reg_acc = reg_o; o0_X = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_73 =>
            -- reg_a = a2_X; reg_b = b5_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_74 =>
            -- reg_a = o2_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_75 =>
            -- reg_a = a3_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_76 =>
            -- reg_a = o3_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_77 =>
            -- reg_a = a4_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_78 =>
            -- reg_a = o4_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_79 =>
            -- reg_a = a5_X; reg_b = b2_X; reg_acc = reg_o; Enable sign a; o1_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_80 =>
            -- reg_a = a3_X; reg_b = b5_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_81 =>
            -- reg_a = o3_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_82 =>
            -- reg_a = a4_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_83 =>
            -- reg_a = o4_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_84 =>
            -- reg_a = a5_X; reg_b = b3_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_85 =>
            -- reg_a = o5_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_86 =>
            -- reg_a = a4_X; reg_b = b5_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_87 =>
            -- reg_a = o4_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_88 =>
            -- reg_a = a5_X; reg_b = b4_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_89 =>
            -- reg_a = o5_X; reg_b = primeSP4; reg_acc = reg_o; o3_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_90 =>
            -- reg_a = a5_X; reg_b = b5_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_91 =>
            -- reg_a = o5_X; reg_b = primeSP5; reg_acc = reg_o; o4_X = reg_o; o5_X = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_93 =>
            -- -- In case of sizes 7, 8
            -- reg_a = a0_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_94 =>
            -- reg_a = a5_X; reg_b = b0_X; reg_acc = reg_o; o5_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_95 =>
            -- reg_a = o0_X; reg_b = primeSP6; reg_acc = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_96 =>
            -- reg_a = a1_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_97 =>
            -- reg_a = o1_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_98 =>
            -- reg_a = a2_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_99 =>
            -- reg_a = o2_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_100 =>
            -- reg_a = a3_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_101 =>
            -- reg_a = o3_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_102 =>
            -- reg_a = a4_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_103 =>
            -- reg_a = a5_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_104 =>
            -- -- In case of size 7
            -- reg_a = a0_X; reg_b = b6_X; reg_acc = reg_o; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_105 =>
            -- reg_a = a6_X; reg_b = b0_X; reg_acc = reg_o; o6_X = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_106 =>
            -- reg_a = a1_X; reg_b = b6_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_107 =>
            -- reg_a = o1_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_108 =>
            -- reg_a = a2_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_109 =>
            -- reg_a = o2_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_110 =>
            -- reg_a = a3_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_111 =>
            -- reg_a = o3_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_112 =>
            -- reg_a = a4_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_113 =>
            -- reg_a = o4_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_114 =>
            -- reg_a = a5_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_115 =>
            -- reg_a = a6_X; reg_b = b1_X; reg_acc = reg_o; o0_X = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_116 =>
            -- reg_a = a2_X; reg_b = b6_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_117 =>
            -- reg_a = o2_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_118 =>
            -- reg_a = a3_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_119 =>
            -- reg_a = o3_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_120 =>
            -- reg_a = a4_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_121 =>
            -- reg_a = o4_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_122 =>
            -- reg_a = a5_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_123 =>
            -- reg_a = o5_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_124 =>
            -- reg_a = a6_X; reg_b = b2_X; reg_acc = reg_o; o1_X = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_125 =>
            -- reg_a = a3_X; reg_b = b6_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_126 =>
            -- reg_a = o3_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_127 =>
            -- reg_a = a4_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_128 =>
            -- reg_a = o4_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_129 =>
            -- reg_a = a5_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_130 =>
            -- reg_a = o5_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_131 =>
            -- reg_a = a6_X; reg_b = b3_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_132 =>
            -- reg_a = o6_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_133 =>
            -- reg_a = a4_X; reg_b = b6_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_134 =>
            -- reg_a = o4_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_135 =>
            -- reg_a = a5_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_136 =>
            -- reg_a = o5_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_137 =>
            -- reg_a = a6_X; reg_b = b4_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_138 =>
            -- reg_a = o6_X; reg_b = primeSP4; reg_acc = reg_o; o3_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_139 =>
            -- reg_a = a5_X; reg_b = b6_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_140 =>
            -- reg_a = o5_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_141 =>
            -- reg_a = a6_X; reg_b = b5_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_142 =>
            -- reg_a = o6_X; reg_b = primeSP5; reg_acc = reg_o; o4_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_143 =>
            -- reg_a = a6_X; reg_b = b6_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_144 =>
            -- reg_a = o6_X; reg_b = primeSP6; reg_acc = reg_o; o5_X = reg_o; o6_X = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_146 =>
            -- -- In case of size 8
            -- reg_a = a0_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_147 =>
            -- reg_a = a6_X; reg_b = b0_X; reg_acc = reg_o; o6_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_148 =>
            -- reg_a = o0_X; reg_b = primeSP7; reg_acc = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_149 =>
            -- reg_a = a1_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_150 =>
            -- reg_a = o1_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_151 =>
            -- reg_a = a2_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_152 =>
            -- reg_a = o2_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_153 =>
            -- reg_a = a3_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_154 =>
            -- reg_a = o3_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_155 =>
            -- reg_a = a4_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_156 =>
            -- reg_a = o4_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_157 =>
            -- reg_a = a5_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_158 =>
            -- reg_a = a6_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_159 =>
            -- reg_a = a0_X; reg_b = b7_X; reg_acc = reg_o; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_160 =>
            -- reg_a = a7_X; reg_b = b0_X; reg_acc = reg_o; o7_X = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "111";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_161 =>
            -- reg_a = a1_X; reg_b = b7_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_162 =>
            -- reg_a = o1_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_163 =>
            -- reg_a = a2_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_164 =>
            -- reg_a = o2_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_165 =>
            -- reg_a = a3_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_166 =>
            -- reg_a = o3_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_167 =>
            -- reg_a = a4_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_168 =>
            -- reg_a = o4_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_169 =>
            -- reg_a = a5_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_170 =>
            -- reg_a = o5_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_171 =>
            -- reg_a = a6_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_172 =>
            -- reg_a = a7_X; reg_b = b1_X; reg_acc = reg_o; o0_X = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_173 =>
            -- reg_a = a2_X; reg_b = b7_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_174 =>
            -- reg_a = o2_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_175 =>
            -- reg_a = a3_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_176 =>
            -- reg_a = o3_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_177 =>
            -- reg_a = a4_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_178 =>
            -- reg_a = o4_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_179 =>
            -- reg_a = a5_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_180 =>
            -- reg_a = o5_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_181 =>
            -- reg_a = a6_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_182 =>
            -- reg_a = o6_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_183 =>
            -- reg_a = a7_X; reg_b = b2_X; reg_acc = reg_o; o1_X = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_184 =>
            -- reg_a = a3_X; reg_b = b7_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_185 =>
            -- reg_a = o3_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_186 =>
            -- reg_a = a4_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_187 =>
            -- reg_a = o4_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_188 =>
            -- reg_a = a5_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_189 =>
            -- reg_a = o5_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_190 =>
            -- reg_a = a6_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_191 =>
            -- reg_a = o6_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_192 =>
            -- reg_a = a7_X; reg_b = b3_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_193 =>
            -- reg_a = o7_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_194 =>
            -- reg_a = a4_X; reg_b = b7_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_195 =>
            -- reg_a = o4_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_196 =>
            -- reg_a = a5_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_197 =>
            -- reg_a = o5_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_198 =>
            -- reg_a = a6_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_199 =>
            -- reg_a = o6_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_200 =>
            -- reg_a = a7_X; reg_b = b4_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_201 =>
            -- reg_a = o7_X; reg_b = primeSP4; reg_acc = reg_o; o3_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_202 =>
            -- reg_a = a5_X; reg_b = b7_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_203 =>
            -- reg_a = o5_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_204 =>
            -- reg_a = a6_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_205 =>
            -- reg_a = o6_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_206 =>
            -- reg_a = a7_X; reg_b = b5_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_207 =>
            -- reg_a = o7_X; reg_b = primeSP5; reg_acc = reg_o; o4_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_208 =>
            -- reg_a = a6_X; reg_b = b7_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_209 =>
            -- reg_a = o6_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_210 =>
            -- reg_a = a7_X; reg_b = b6_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_211 =>
            -- reg_a = o7_X; reg_b = primeSP6; reg_acc = reg_o; o5_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_212 =>
            -- reg_a = a7_X; reg_b = b7_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_213 =>
            -- reg_a = o7_X; reg_b = primeSP7; reg_acc = reg_o; o6_X = reg_o; o7_X = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_0 =>
            -- -- In case of size 1
            -- reg_a = a0_X; reg_b = a0_X; reg_acc = 0; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_1 =>
            -- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o0_X = reg_y; operation : keep accumulator;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "11";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "10";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "11";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '1';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_2 =>
            -- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "01";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_3 =>
            -- reg_a = 0; reg_b = 0; reg_acc = reg_o >> 256; o0_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "11";
            next_mac_clear_reg_b <= '1';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_5 =>
            -- -- In case of 2, 3, 4, 5, 6, 7, 8
            -- reg_a = a0_X; reg_b = a0_X; reg_acc = 0; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_6 =>
            -- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o0_X = reg_y; operation : keep accumulator;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "11";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "10";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "11";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '1';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_7 =>
            -- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "01";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_8 =>
            -- reg_a = o0_X; reg_b = prime1; reg_acc = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_9 =>
            -- -- In case of size 2
            -- reg_a = a0_X; reg_b = a1_X; reg_acc = reg_o; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_10 =>
            -- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o1_X = reg_y; operation : keep accumulator;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "11";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "10";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "11";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '1';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_11 =>
            -- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "01";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_12 =>
            -- reg_a = a1_X; reg_b = a1_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_13 =>
            -- reg_a = o1_X; reg_b = prime1; reg_acc = reg_o; o0_X = reg_o; o1_X = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_15 =>
            -- -- Others cases
            -- reg_a = a0_X; reg_b = a1_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_16 =>
            -- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o1_X = reg_y; operation : keep accumulator;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "11";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "10";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "11";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '1';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_17 =>
            -- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "01";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_18 =>
            -- reg_a = o0_X; reg_b = prime2; reg_acc = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_19 =>
            -- reg_a = a1_X; reg_b = a1_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_20 =>
            -- reg_a = o1_X; reg_b = prime1; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_21 =>
            -- -- In case of size 3
            -- reg_a = a0_X; reg_b = a2_X; reg_acc = reg_o; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_22 =>
            -- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o2_X = reg_y; operation : keep accumulator;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "11";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "10";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "11";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '1';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_23 =>
            -- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "01";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_24 =>
            -- reg_a = a1_X; reg_b = a2_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_25 =>
            -- reg_a = o1_X; reg_b = prime2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_26 =>
            -- reg_a = o2_X; reg_b = prime1; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_27 =>
            -- reg_a = a2_X; reg_b = a2_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_28 =>
            -- reg_a = o2_X; reg_b = prime2; reg_acc = reg_o; o1_X = reg_o; o2_X = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_30 =>
            -- -- Other cases
            -- reg_a = a0_X; reg_b = a2_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_31 =>
            -- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o2_X = reg_y; operation : keep accumulator;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "11";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "10";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "11";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '1';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_32 =>
            -- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "01";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_33 =>
            -- reg_a = o0_X; reg_b = prime3; reg_acc = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_34 =>
            -- reg_a = a1_X; reg_b = a2_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_35 =>
            -- reg_a = o1_X; reg_b = prime2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_36 =>
            -- reg_a = o2_X; reg_b = prime1; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_37 =>
            -- In case of size 4
            -- reg_a = a0_X; reg_b = a3_X; reg_acc = reg_o; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_38 =>
            -- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o3_X = reg_y; operation : keep accumulator;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "11";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "10";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "11";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '1';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_39 =>
            -- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "01";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_40 =>
            -- reg_a = a1_X; reg_b = a3_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_41 =>
            -- reg_a = o1_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_42 =>
            -- reg_a = a2_X; reg_b = a2_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_43 =>
            -- reg_a = o2_X; reg_b = prime2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_44 =>
            -- reg_a = o3_X; reg_b = prime1; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_45 =>
            -- reg_a = a2_X; reg_b = a3_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_46 =>
            -- reg_a = o2_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_47 =>
            -- reg_a = o3_X; reg_b = prime2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_48 =>
            -- reg_a = a3_X; reg_b = a3_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_49 =>
            -- reg_a = o3_X; reg_b = prime3; reg_acc = reg_o; o2_X = reg_o; o3_X = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_51 =>
            -- -- Other cases
            -- reg_a = a0_X; reg_b = a3_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_52 =>
            -- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o3_X = reg_y; operation : keep accumulator;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "11";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "10";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "11";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '1';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_53 =>
            -- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "01";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_54 =>
            -- reg_a = o0_X; reg_b = prime4; reg_acc = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_55 =>
            -- reg_a = a1_X; reg_b = a3_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_56 =>
            -- reg_a = o1_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_57 =>
            -- reg_a = a2_X; reg_b = a2_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_58 =>
            -- reg_a = o2_X; reg_b = prime2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_59 =>
            -- reg_a = o3_X; reg_b = prime1; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_60 =>
            -- -- In case of size 5
            -- reg_a = a0_X; reg_b = a4_X; reg_acc = reg_o; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_61 =>
            -- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o4_X = reg_y; operation : keep accumulator;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "11";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "10";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "11";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '1';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_62 =>
            -- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "01";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_63 =>
            -- reg_a = a1_X; reg_b = a4_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_64 =>
            -- reg_a = o1_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_65 =>
            -- reg_a = a2_X; reg_b = a3_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_66 =>
            -- reg_a = o2_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_67 =>
            -- reg_a = o3_X; reg_b = prime2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_68 =>
            -- reg_a = o4_X; reg_b = prime1; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_69 =>
            -- reg_a = a2_X; reg_b = a4_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_70 =>
            -- reg_a = o2_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_71 =>
            -- reg_a = a3_X; reg_b = a3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_72 =>
            -- reg_a = o3_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_73 =>
            -- reg_a = o4_X; reg_b = prime2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_74 =>
            -- reg_a = a3_X; reg_b = a4_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_75 =>
            -- reg_a = o3_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_76 =>
            -- reg_a = o4_X; reg_b = prime3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_77 =>
            -- reg_a = a4_X; reg_b = a4_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_78 =>
            -- reg_a = o4_X; reg_b = prime4; reg_acc = reg_o; o3_X = reg_o; o4_X = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_80 =>
            -- -- Other cases
            -- reg_a = a0_X; reg_b = a4_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_81 =>
            -- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o4_X = reg_y; operation : keep accumulator;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "11";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "10";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "11";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '1';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_82 =>
            -- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "01";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_83 =>
            -- reg_a = o0_X; reg_b = prime5; reg_acc = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_84 =>
            -- reg_a = a1_X; reg_b = a4_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_85 =>
            -- reg_a = o1_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_86 =>
            -- reg_a = a2_X; reg_b = a3_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_87 =>
            -- reg_a = o2_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_88 =>
            -- reg_a = o3_X; reg_b = prime2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_89 =>
            -- reg_a = o4_X; reg_b = prime1; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_90 =>
            -- -- In case of size 6
            -- reg_a = a0_X; reg_b = a5_X; reg_acc = reg_o; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_91 =>
            -- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o5_X = reg_y; operation : keep accumulator;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "11";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "10";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "11";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '1';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_92 =>
            -- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "01";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_93 =>
            -- reg_a = a1_X; reg_b = a5_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_94 =>
            -- reg_a = o1_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_95 =>
            -- reg_a = a2_X; reg_b = a4_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_96 =>
            -- reg_a = o2_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_97 =>
            -- reg_a = a3_X; reg_b = a3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_98 =>
            -- reg_a = o3_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_99 =>
            -- reg_a = o4_X; reg_b = prime2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_100 =>
            -- reg_a = o5_X; reg_b = prime1; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_101 =>
            -- reg_a = a2_X; reg_b = a5_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_102 =>
            -- reg_a = o2_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_103 =>
            -- reg_a = a3_X; reg_b = a4_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_104 =>
            -- reg_a = o3_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_105 =>
            -- reg_a = o4_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_106 =>
            -- reg_a = o5_X; reg_b = prime2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_107 =>
            -- reg_a = a3_X; reg_b = a5_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_108 =>
            -- reg_a = o3_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_109 =>
            -- reg_a = a4_X; reg_b = a4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_110 =>
            -- reg_a = o4_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_111 =>
            -- reg_a = o5_X; reg_b = prime3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_112 =>
            -- reg_a = a4_X; reg_b = a5_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_113 =>
            -- reg_a = o4_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_114 =>
            -- reg_a = o5_X; reg_b = prime4; reg_acc = reg_o; o3_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_115 =>
            -- reg_a = a5_X; reg_b = a5_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_116 =>
            -- reg_a = o5_X; reg_b = prime5; reg_acc = reg_o; o4_X = reg_o; o5_X = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_118 =>
            -- -- Other cases
            -- reg_a = a0_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_119 =>
            -- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o5_X = reg_y; operation : keep accumulator;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "11";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "10";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "11";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '1';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_120 =>
            -- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "01";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_121 =>
            -- reg_a = o0_X; reg_b = prime6; reg_acc = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_122 =>
            -- reg_a = a1_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_123 =>
            -- reg_a = o1_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_124 =>
            -- reg_a = a2_X; reg_b = a4_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_125 =>
            -- reg_a = o2_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_126 =>
            -- reg_a = a3_X; reg_b = a3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_127 =>
            -- reg_a = o3_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_128 =>
            -- reg_a = o4_X; reg_b = prime2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_129 =>
            -- reg_a = o5_X; reg_b = prime1; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_130 =>
            -- -- In case of size 7
            -- reg_a = a0_X; reg_b = a6_X; reg_acc = reg_o; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_131 =>
            -- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o6_X = reg_y; operation : keep accumulator;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "11";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "10";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "11";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '1';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_132 =>
            -- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "01";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_133 =>
            -- reg_a = a1_X; reg_b = a6_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_134 =>
            -- reg_a = o1_X; reg_b = prime6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_135 =>
            -- reg_a = a2_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_136 =>
            -- reg_a = o2_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_137 =>
            -- reg_a = a3_X; reg_b = a4_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_138 =>
            -- reg_a = o3_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_139 =>
            -- reg_a = o4_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_140 =>
            -- reg_a = o5_X; reg_b = prime2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_141 =>
            -- reg_a = o6_X; reg_b = prime1; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_142 =>
            -- reg_a = a2_X; reg_b = a6_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_143 =>
            -- reg_a = o2_X; reg_b = prime6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_144 =>
            -- reg_a = a3_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_145 =>
            -- reg_a = o3_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_146 =>
            -- reg_a = a4_X; reg_b = a4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_147 =>
            -- reg_a = o4_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_148 =>
            -- reg_a = o5_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_149 =>
            -- reg_a = o6_X; reg_b = prime2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_150 =>
            -- reg_a = a3_X; reg_b = a6_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_151 =>
            -- reg_a = o3_X; reg_b = prime6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_152 =>
            -- reg_a = a4_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_153 =>
            -- reg_a = o4_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_154 =>
            -- reg_a = o5_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_155 =>
            -- reg_a = o6_X; reg_b = prime3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_156 =>
            -- reg_a = a4_X; reg_b = a6_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_157 =>
            -- reg_a = o4_X; reg_b = prime6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_158 =>
            -- reg_a = a5_X; reg_b = a5_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_159 =>
            -- reg_a = o5_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_160 =>
            -- reg_a = o6_X; reg_b = prime4; reg_acc = reg_o; o3_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_161 =>
            -- reg_a = a5_X; reg_b = a6_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_162 =>
            -- reg_a = o5_X; reg_b = prime6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_163 =>
            -- reg_a = o6_X; reg_b = prime5; reg_acc = reg_o; o4_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_164 =>
            -- reg_a = a6_X; reg_b = a6_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_165 =>
            -- reg_a = o6_X; reg_b = prime6; reg_acc = reg_o; o5_X = reg_o; o6_X = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_167 =>
            -- -- In case of size 8
            -- reg_a = a0_X; reg_b = a6_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_168 =>
            -- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o6_X = reg_y; operation : keep accumulator;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "11";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "10";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "11";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '1';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_169 =>
            -- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "01";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_170 =>
            -- reg_a = o0_X; reg_b = prime7; reg_acc = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_171 =>
            -- reg_a = a1_X; reg_b = a6_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_172 =>
            -- reg_a = o1_X; reg_b = prime6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_173 =>
            -- reg_a = a2_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_174 =>
            -- reg_a = o2_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_175 =>
            -- reg_a = a3_X; reg_b = a4_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_176 =>
            -- reg_a = o3_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_177 =>
            -- reg_a = o4_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_178 =>
            -- reg_a = o5_X; reg_b = prime2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_179 =>
            -- reg_a = o6_X; reg_b = prime1; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_180 =>
            -- reg_a = a0_X; reg_b = a7_X; reg_acc = reg_o; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_181 =>
            -- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o7_X = reg_y; operation : keep accumulator;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "11";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "111";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "10";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "11";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '1';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_182 =>
            -- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "01";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_183 =>
            -- reg_a = a1_X; reg_b = a7_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_184 =>
            -- reg_a = o1_X; reg_b = prime7; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_185 =>
            -- reg_a = a2_X; reg_b = a6_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_186 =>
            -- reg_a = o2_X; reg_b = prime6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_187 =>
            -- reg_a = a3_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_188 =>
            -- reg_a = o3_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_189 =>
            -- reg_a = a4_X; reg_b = a4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_190 =>
            -- reg_a = o4_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_191 =>
            -- reg_a = o5_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_192 =>
            -- reg_a = o6_X; reg_b = prime2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_193 =>
            -- reg_a = o7_X; reg_b = prime1; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_194 =>
            -- reg_a = a2_X; reg_b = a7_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_195 =>
            -- reg_a = o2_X; reg_b = prime7; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_196 =>
            -- reg_a = a3_X; reg_b = a6_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_197 =>
            -- reg_a = o3_X; reg_b = prime6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_198 =>
            -- reg_a = a4_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_199 =>
            -- reg_a = o4_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_200 =>
            -- reg_a = o5_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_201 =>
            -- reg_a = o6_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_202 =>
            -- reg_a = o7_X; reg_b = prime2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_203 =>
            -- reg_a = a3_X; reg_b = a7_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_204 =>
            -- reg_a = o3_X; reg_b = prime7; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_205 =>
            -- reg_a = a4_X; reg_b = a6_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_206 =>
            -- reg_a = o4_X; reg_b = prime6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_207 =>
            -- reg_a = a5_X; reg_b = a5_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_208 =>
            -- reg_a = o5_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_209 =>
            -- reg_a = o6_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_210 =>
            -- reg_a = o7_X; reg_b = prime3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_211 =>
            -- reg_a = a4_X; reg_b = a7_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_212 =>
            -- reg_a = o4_X; reg_b = prime7; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_213 =>
            -- reg_a = a5_X; reg_b = a6_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_214 =>
            -- reg_a = o5_X; reg_b = prime6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_215 =>
            -- reg_a = o6_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_216 =>
            -- reg_a = o7_X; reg_b = prime4; reg_acc = reg_o; o3_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_217 =>
            -- reg_a = a5_X; reg_b = a7_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_218 =>
            -- reg_a = o5_X; reg_b = prime7; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_219 =>
            -- reg_a = a6_X; reg_b = a6_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_220 =>
            -- reg_a = o6_X; reg_b = prime6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_221 =>
            -- reg_a = o7_X; reg_b = prime5; reg_acc = reg_o; o4_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_222 =>
            -- reg_a = a6_X; reg_b = a7_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_223 =>
            -- reg_a = o6_X; reg_b = prime7; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_224 =>
            -- reg_a = o7_X; reg_b = prime6; reg_acc = reg_o; o5_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_225 =>
            -- reg_a = a7_X; reg_b = a7_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_226 =>
            -- reg_a = o7_X; reg_b = prime7; reg_acc = reg_o; o6_X = reg_o; o7_X = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_0 =>
            -- -- In case of size 1
            -- reg_a = a0_X; reg_b = a0_X; reg_acc = 0; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_1 =>
            -- reg_a = 0; reg_b = 0; reg_acc = reg_o >> 256; o0_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "11";
            next_mac_clear_reg_b <= '1';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_3 =>
            -- -- In case of size 2, 3, 4, 5, 6, 7, 8
            -- reg_a = a0_X; reg_b = a0_X; reg_acc = 0; o0_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_4 =>
            -- reg_a = reg_o; reg_b = primeSP1; reg_acc = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "10";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_5 =>
            -- -- In case of size 2
            -- reg_a = a0_X; reg_b = a1_X; reg_acc = reg_o; o1_X = reg_o; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_6 =>
            -- reg_a = a1_X; reg_b = a1_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_7 =>
            -- reg_a = o1_X; reg_b = primeSP1; reg_acc = reg_o; o0_X = reg_o; o1_X = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_9 =>
            -- -- In case of size 3, 4, 5, 6, 7, 8
            -- reg_a = a0_X; reg_b = a1_X; reg_acc = reg_o; o1_X = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_10 =>
            -- reg_a = o0_X; reg_b = primeSP2; reg_acc = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_11 =>
            -- reg_a = a1_X; reg_b = a1_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_12 =>
            -- reg_a = o1_X; reg_b = primeSP1; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_13 =>
            -- -- In case of size 3
            -- reg_a = a0_X; reg_b = a2_X; reg_acc = reg_o; o2_X = reg_o; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_14 =>
            -- reg_a = a1_X; reg_b = a2_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_15 =>
            -- reg_a = o1_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_16 =>
            -- reg_a = o2_X; reg_b = primeSP1; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_17 =>
            -- reg_a = a2_X; reg_b = a2_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_18 =>
            -- reg_a = o2_X; reg_b = primeSP2; reg_acc = reg_o; o1_X = reg_o; o2_X = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_20 =>
            -- -- In case of sizes 4, 5, 6, 7, 8
            -- reg_a = a0_X; reg_b = a2_X; reg_acc = reg_o; o2_X = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_21 =>
            -- reg_a = o0_X; reg_b = primeSP3; reg_acc = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_22 =>
            -- reg_a = a1_X; reg_b = a2_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_23 =>
            -- reg_a = o1_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_24 =>
            -- reg_a = o2_X; reg_b = primeSP1; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_25 =>
            -- -- In case of size 4
            -- reg_a = a0_X; reg_b = a3_X; reg_acc = reg_o; o3_X = reg_o; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_26 =>
            -- reg_a = a1_X; reg_b = a3_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_27 =>
            -- reg_a = o1_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_28 =>
            -- reg_a = a2_X; reg_b = a2_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_29 =>
            -- reg_a = o2_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_30 =>
            -- reg_a = o3_X; reg_b = primeSP1; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_31 =>
            -- reg_a = a2_X; reg_b = a3_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_32 =>
            -- reg_a = o2_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_33 =>
            -- reg_a = o3_X; reg_b = primeSP2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_34 =>
            -- reg_a = a3_X; reg_b = a3_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_35 =>
            -- reg_a = o3_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; o3_X = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_37 =>
            -- -- In case of sizes 5, 6, 7, 8
            -- reg_a = a0_X; reg_b = a3_X; reg_acc = reg_o; o3_X = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_38 =>
            -- reg_a = o0_X; reg_b = primeSP4; reg_acc = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_39 =>
            -- reg_a = a1_X; reg_b = a3_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_40 =>
            -- reg_a = o1_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_41 =>
            -- reg_a = a2_X; reg_b = a2_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_42 =>
            -- reg_a = o2_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_43 =>
            -- reg_a = o3_X; reg_b = primeSP1; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_44 =>
            -- -- In case of size 5
            -- reg_a = a0_X; reg_b = a4_X; reg_acc = reg_o; o4_X = reg_o; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_45 =>
            -- reg_a = a1_X; reg_b = a4_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_46 =>
            -- reg_a = o1_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_47 =>
            -- reg_a = a2_X; reg_b = a3_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_48 =>
            -- reg_a = o2_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_49 =>
            -- reg_a = o3_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_50 =>
            -- reg_a = o4_X; reg_b = primeSP1; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_51 =>
            -- reg_a = a2_X; reg_b = a4_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_52 =>
            -- reg_a = o2_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_53 =>
            -- reg_a = a3_X; reg_b = a3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_54 =>
            -- reg_a = o3_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_55 =>
            -- reg_a = o4_X; reg_b = primeSP2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_56 =>
            -- reg_a = a3_X; reg_b = a4_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_57 =>
            -- reg_a = o3_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_58 =>
            -- reg_a = o4_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_59 =>
            -- reg_a = a4_X; reg_b = a4_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_60 =>
            -- reg_a = o4_X; reg_b = primeSP4; reg_acc = reg_o; o3_X = reg_o; o4_X = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_62 =>
            -- -- In case of sizes 6, 7, 8
            -- reg_a = a0_X; reg_b = a4_X; reg_acc = reg_o; o4_X = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_63 =>
            -- reg_a = o0_X; reg_b = primeSP5; reg_acc = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_64 =>
            -- reg_a = a1_X; reg_b = a4_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_65 =>
            -- reg_a = o1_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_66 =>
            -- reg_a = a2_X; reg_b = a3_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_67 =>
            -- reg_a = o2_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_68 =>
            -- reg_a = o3_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_69 =>
            -- reg_a = o4_X; reg_b = primeSP1; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_70 =>
            -- -- In case of size 6
            -- reg_a = a0_X; reg_b = a5_X; reg_acc = reg_o; o5_X = reg_o; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_71 =>
            -- reg_a = a1_X; reg_b = a5_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_72 =>
            -- reg_a = o1_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_73 =>
            -- reg_a = a2_X; reg_b = a4_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_74 =>
            -- reg_a = o2_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_75 =>
            -- reg_a = a3_X; reg_b = a3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_76 =>
            -- reg_a = o3_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_77 =>
            -- reg_a = o4_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_78 =>
            -- reg_a = o5_X; reg_b = primeSP1; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_79 =>
            -- reg_a = a2_X; reg_b = a5_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_80 =>
            -- reg_a = o2_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_81 =>
            -- reg_a = a3_X; reg_b = a4_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_82 =>
            -- reg_a = o3_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_83 =>
            -- reg_a = o4_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_84 =>
            -- reg_a = o5_X; reg_b = primeSP2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_85 =>
            -- reg_a = a3_X; reg_b = a5_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_86 =>
            -- reg_a = o3_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_87 =>
            -- reg_a = a4_X; reg_b = a4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_88 =>
            -- reg_a = o4_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_89 =>
            -- reg_a = o5_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_90 =>
            -- reg_a = a4_X; reg_b = a5_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_91 =>
            -- reg_a = o4_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_92 =>
            -- reg_a = o5_X; reg_b = primeSP4; reg_acc = reg_o; o3_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_93 =>
            -- reg_a = a5_X; reg_b = a5_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_94 =>
            -- reg_a = o5_X; reg_b = primeSP5; reg_acc = reg_o; o4_X = reg_o; o5_X = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_96 =>
            -- -- In case of sizes 7, 8
            -- reg_a = a0_X; reg_b = a5_X; reg_acc = reg_o; o5_X = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_97 =>
            -- reg_a = o0_X; reg_b = primeSP6; reg_acc = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_98 =>
            -- reg_a = a1_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_99 =>
            -- reg_a = o1_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_100 =>
            -- reg_a = a2_X; reg_b = a4_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_101 =>
            -- reg_a = o2_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_102 =>
            -- reg_a = a3_X; reg_b = a3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_103 =>
            -- reg_a = o3_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_104 =>
            -- reg_a = o4_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_105 =>
            -- reg_a = o5_X; reg_b = primeSP1; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_106 =>
            -- -- In case of size 7
            -- reg_a = a0_X; reg_b = a6_X; reg_acc = reg_o; o6_X = reg_o; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_107 =>
            -- reg_a = a1_X; reg_b = a6_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_108 =>
            -- reg_a = o1_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_109 =>
            -- reg_a = a2_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_110 =>
            -- reg_a = o2_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_111 =>
            -- reg_a = a3_X; reg_b = a4_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_112 =>
            -- reg_a = o3_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_113 =>
            -- reg_a = o4_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_114 =>
            -- reg_a = o5_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_115 =>
            -- reg_a = o6_X; reg_b = primeSP1; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_116 =>
            -- reg_a = a2_X; reg_b = a6_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_117 =>
            -- reg_a = o2_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_118 =>
            -- reg_a = a3_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_119 =>
            -- reg_a = o3_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_120 =>
            -- reg_a = a4_X; reg_b = a4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_121 =>
            -- reg_a = o4_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_122 =>
            -- reg_a = o5_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_123 =>
            -- reg_a = o6_X; reg_b = primeSP2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_124 =>
            -- reg_a = a3_X; reg_b = a6_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_125 =>
            -- reg_a = o3_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_126 =>
            -- reg_a = a4_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_127 =>
            -- reg_a = o4_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_128 =>
            -- reg_a = o5_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_129 =>
            -- reg_a = o6_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_130 =>
            -- reg_a = a4_X; reg_b = a6_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_131 =>
            -- reg_a = o4_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_132 =>
            -- reg_a = a5_X; reg_b = a5_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_133 =>
            -- reg_a = o5_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_134 =>
            -- reg_a = o6_X; reg_b = primeSP4; reg_acc = reg_o; o3_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_135 =>
            -- reg_a = a5_X; reg_b = a6_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_136 =>
            -- reg_a = o5_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_137 =>
            -- reg_a = o6_X; reg_b = primeSP5; reg_acc = reg_o; o4_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_138 =>
            -- reg_a = a6_X; reg_b = a6_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_139 =>
            -- reg_a = o6_X; reg_b = primeSP6; reg_acc = reg_o; o5_X = reg_o; o6_X = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_141 =>
            -- -- In case of size 8
            -- reg_a = a0_X; reg_b = a6_X; reg_acc = reg_o; o6_X = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_142 =>
            -- reg_a = o0_X; reg_b = primeSP7; reg_acc = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_143 =>
            -- reg_a = a1_X; reg_b = a6_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_144 =>
            -- reg_a = o1_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_145 =>
            -- reg_a = a2_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_146 =>
            -- reg_a = o2_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_147 =>
            -- reg_a = a3_X; reg_b = a4_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_148 =>
            -- reg_a = o3_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_149 =>
            -- reg_a = o4_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_150 =>
            -- reg_a = o5_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_151 =>
            -- reg_a = o6_X; reg_b = primeSP1; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_152 =>
            -- reg_a = a0_X; reg_b = a7_X; reg_acc = reg_o; o7_X = reg_o; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "111";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_153 =>
            -- reg_a = a1_X; reg_b = a7_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_154 =>
            -- reg_a = o1_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_155 =>
            -- reg_a = a2_X; reg_b = a6_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_156 =>
            -- reg_a = o2_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_157 =>
            -- reg_a = a3_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_158 =>
            -- reg_a = o3_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_159 =>
            -- reg_a = a4_X; reg_b = a4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_160 =>
            -- reg_a = o4_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_161 =>
            -- reg_a = o5_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_162 =>
            -- reg_a = o6_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_163 =>
            -- reg_a = o7_X; reg_b = primeSP1; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_164 =>
            -- reg_a = a2_X; reg_b = a7_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_165 =>
            -- reg_a = o2_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_166 =>
            -- reg_a = a3_X; reg_b = a6_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_167 =>
            -- reg_a = o3_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_168 =>
            -- reg_a = a4_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_169 =>
            -- reg_a = o4_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_170 =>
            -- reg_a = o5_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_171 =>
            -- reg_a = o6_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_172 =>
            -- reg_a = o7_X; reg_b = primeSP2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_173 =>
            -- reg_a = a3_X; reg_b = a7_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_174 =>
            -- reg_a = o3_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_175 =>
            -- reg_a = a4_X; reg_b = a6_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_176 =>
            -- reg_a = o4_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_177 =>
            -- reg_a = a5_X; reg_b = a5_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_178 =>
            -- reg_a = o5_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_179 =>
            -- reg_a = o6_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_180 =>
            -- reg_a = o7_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_181 =>
            -- reg_a = a4_X; reg_b = a7_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_182 =>
            -- reg_a = o4_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_183 =>
            -- reg_a = a5_X; reg_b = a6_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_184 =>
            -- reg_a = o5_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_185 =>
            -- reg_a = o6_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_186 =>
            -- reg_a = o7_X; reg_b = primeSP4; reg_acc = reg_o; o3_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_187 =>
            -- reg_a = a5_X; reg_b = a7_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_188 =>
            -- reg_a = o5_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_189 =>
            -- reg_a = a6_X; reg_b = a6_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_190 =>
            -- reg_a = o6_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_191 =>
            -- reg_a = o7_X; reg_b = primeSP5; reg_acc = reg_o; o4_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_192 =>
            -- reg_a = a6_X; reg_b = a7_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_193 =>
            -- reg_a = o6_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_194 =>
            -- reg_a = o7_X; reg_b = primeSP6; reg_acc = reg_o; o5_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_195 =>
            -- reg_a = a7_X; reg_b = a7_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_196 =>
            -- reg_a = o7_X; reg_b = primeSP7; reg_acc = reg_o; o6_X = reg_o; o7_X = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_0 =>
            -- -- In case of size 2, 3, 4, 5, 6, 7, 8
            -- reg_a = a0_X; reg_b = a0_X; reg_acc = 0; o0_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_1 =>
            -- -- In case of size 2
            -- reg_a = a0_X; reg_b = a1_X; reg_acc = reg_o; o1_X = reg_o; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_2 =>
            -- reg_a = a1_X; reg_b = a1_X; reg_acc = reg_o >> 256; Enable sign a,b; o0_X = reg_o; o1_X = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_4 =>
            -- -- In case of size 3, 4, 5, 6, 7, 8
            -- reg_a = a0_X; reg_b = a1_X; reg_acc = reg_o >> 256; o1_X = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_5 =>
            -- reg_a = o0_X; reg_b = primeSP2; reg_acc = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_6 =>
            -- reg_a = a1_X; reg_b = a1_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_7 =>
            -- -- In case of size 3
            -- reg_a = a0_X; reg_b = a2_X; reg_acc = reg_o; o2_X = reg_o; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_8 =>
            -- reg_a = a1_X; reg_b = a2_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_9 =>
            -- reg_a = o1_X; reg_b = primeSP2; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_10 =>
            -- reg_a = a2_X; reg_b = a2_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_11 =>
            -- reg_a = o2_X; reg_b = primeSP2; reg_acc = reg_o; o1_X = reg_o; o2_X = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_13 =>
            -- -- In case of size 4, 5, 6, 7, 8
            -- reg_a = a0_X; reg_b = a2_X; reg_acc = reg_o; o2_X = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_14 =>
            -- reg_a = o0_X; reg_b = primeSP3; reg_acc = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_15 =>
            -- reg_a = a1_X; reg_b = a2_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_16 =>
            -- reg_a = o1_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_17 =>
            -- -- In case of size 4
            -- reg_a = a0_X; reg_b = a3_X; reg_acc = reg_o; o3_X = reg_o; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_18 =>
            -- reg_a = a1_X; reg_b = a3_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_19 =>
            -- reg_a = o1_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_20 =>
            -- reg_a = a2_X; reg_b = a2_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_21 =>
            -- reg_a = o2_X; reg_b = primeSP2; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_22 =>
            -- reg_a = a2_X; reg_b = a3_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_23 =>
            -- reg_a = o2_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_24 =>
            -- reg_a = o3_X; reg_b = primeSP2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_25 =>
            -- reg_a = a3_X; reg_b = a3_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_26 =>
            -- reg_a = o3_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; o3_X = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_28 =>
            -- -- In case of size 5, 6, 7, 8
            -- reg_a = a0_X; reg_b = a3_X; reg_acc = reg_o; o3_X = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_29 =>
            -- reg_a = o0_X; reg_b = primeSP4; reg_acc = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_30 =>
            -- reg_a = a1_X; reg_b = a3_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_31 =>
            -- reg_a = o1_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_32 =>
            -- reg_a = a2_X; reg_b = a2_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_33 =>
            -- reg_a = o2_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_34 =>
            -- -- In case of size 5
            -- reg_a = a0_X; reg_b = a4_X; reg_acc = reg_o; o4_X = reg_o; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_35 =>
            -- reg_a = a1_X; reg_b = a4_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_36 =>
            -- reg_a = o1_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_37 =>
            -- reg_a = a2_X; reg_b = a3_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_38 =>
            -- reg_a = o2_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_39 =>
            -- reg_a = o3_X; reg_b = primeSP2; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_40 =>
            -- reg_a = a2_X; reg_b = a4_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_41 =>
            -- reg_a = o2_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_42 =>
            -- reg_a = a3_X; reg_b = a3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_43 =>
            -- reg_a = o3_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_44 =>
            -- reg_a = o4_X; reg_b = primeSP2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_45 =>
            -- reg_a = a3_X; reg_b = a4_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_46 =>
            -- reg_a = o3_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_47 =>
            -- reg_a = o4_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_48 =>
            -- reg_a = a4_X; reg_b = a4_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_49 =>
            -- reg_a = o4_X; reg_b = primeSP4; reg_acc = reg_o; o3_X = reg_o; o4_X = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_51 =>
            -- -- In case of sizes 6, 7, 8
            -- reg_a = a0_X; reg_b = a4_X; reg_acc = reg_o; o4_X = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_52 =>
            -- reg_a = o0_X; reg_b = primeSP5; reg_acc = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_53 =>
            -- reg_a = a1_X; reg_b = a4_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_54 =>
            -- reg_a = o1_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_55 =>
            -- reg_a = a2_X; reg_b = a3_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_56 =>
            -- reg_a = o2_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_57 =>
            -- reg_a = o3_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_58 =>
            -- -- In case of size 6
            -- reg_a = a0_X; reg_b = a5_X; reg_acc = reg_o; o5_X = reg_o; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_59 =>
            -- reg_a = a1_X; reg_b = a5_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_60 =>
            -- reg_a = o1_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_61 =>
            -- reg_a = a2_X; reg_b = a4_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_62 =>
            -- reg_a = o2_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_63 =>
            -- reg_a = a3_X; reg_b = a3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_64 =>
            -- reg_a = o3_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_65 =>
            -- reg_a = o4_X; reg_b = primeSP2; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_66 =>
            -- reg_a = a2_X; reg_b = a5_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_67 =>
            -- reg_a = o2_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_68 =>
            -- reg_a = a3_X; reg_b = a4_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_69 =>
            -- reg_a = o3_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_70 =>
            -- reg_a = o4_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_71 =>
            -- reg_a = o5_X; reg_b = primeSP2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_72 =>
            -- reg_a = a3_X; reg_b = a5_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_73 =>
            -- reg_a = o3_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_74 =>
            -- reg_a = a4_X; reg_b = a4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_75 =>
            -- reg_a = o4_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_76 =>
            -- reg_a = o5_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_77 =>
            -- reg_a = a4_X; reg_b = a5_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_78 =>
            -- reg_a = o4_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_79 =>
            -- reg_a = o5_X; reg_b = primeSP4; reg_acc = reg_o; o3_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_80 =>
            -- reg_a = a5_X; reg_b = a5_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_81 =>
            -- reg_a = o5_X; reg_b = primeSP5; reg_acc = reg_o; o4_X = reg_o; o5_X = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_83 =>
            -- -- In case of sizes 7, 8
            -- reg_a = a0_X; reg_b = a5_X; reg_acc = reg_o; o5_X = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_84 =>
            -- reg_a = o0_X; reg_b = primeSP6; reg_acc = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_85 =>
            -- reg_a = a1_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_86 =>
            -- reg_a = o1_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_87 =>
            -- reg_a = a2_X; reg_b = a4_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_88 =>
            -- reg_a = o2_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_89 =>
            -- reg_a = a3_X; reg_b = a3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_90 =>
            -- reg_a = o3_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_91 =>
            -- reg_a = o4_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_92 =>
            -- -- In case of size 7
            -- reg_a = a0_X; reg_b = a6_X; reg_acc = reg_o; o6_X = reg_o; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_93 =>
            -- reg_a = a1_X; reg_b = a6_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_94 =>
            -- reg_a = o1_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_95 =>
            -- reg_a = a2_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_96 =>
            -- reg_a = o2_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_97 =>
            -- reg_a = a3_X; reg_b = a4_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_98 =>
            -- reg_a = o3_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_99 =>
            -- reg_a = o4_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_100 =>
            -- reg_a = o5_X; reg_b = primeSP2; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_101 =>
            -- reg_a = a2_X; reg_b = a6_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_102 =>
            -- reg_a = o2_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_103 =>
            -- reg_a = a3_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_104 =>
            -- reg_a = o3_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_105 =>
            -- reg_a = a4_X; reg_b = a4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_106 =>
            -- reg_a = o4_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_107 =>
            -- reg_a = o5_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_108 =>
            -- reg_a = o6_X; reg_b = primeSP2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_109 =>
            -- reg_a = a3_X; reg_b = a6_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_110 =>
            -- reg_a = o3_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_111 =>
            -- reg_a = a4_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_112 =>
            -- reg_a = o4_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_113 =>
            -- reg_a = o5_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_114 =>
            -- reg_a = o6_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_115 =>
            -- reg_a = a4_X; reg_b = a6_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_116 =>
            -- reg_a = o4_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_117 =>
            -- reg_a = a5_X; reg_b = a5_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_118 =>
            -- reg_a = o5_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_119 =>
            -- reg_a = o6_X; reg_b = primeSP4; reg_acc = reg_o; o3_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_120 =>
            -- reg_a = a5_X; reg_b = a6_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_121 =>
            -- reg_a = o5_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_122 =>
            -- reg_a = o6_X; reg_b = primeSP5; reg_acc = reg_o; o4_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_123 =>
            -- reg_a = a6_X; reg_b = a6_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_124 =>
            -- reg_a = o6_X; reg_b = primeSP6; reg_acc = reg_o; o5_X = reg_o; o6_X = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_126 =>
            -- -- In case of size 8
            -- reg_a = a0_X; reg_b = a6_X; reg_acc = reg_o; o6_X = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_127 =>
            -- reg_a = o0_X; reg_b = primeSP7; reg_acc = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_128 =>
            -- reg_a = a1_X; reg_b = a6_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_129 =>
            -- reg_a = o1_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_130 =>
            -- reg_a = a2_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_131 =>
            -- reg_a = o2_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_132 =>
            -- reg_a = a3_X; reg_b = a4_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_133 =>
            -- reg_a = o3_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_134 =>
            -- reg_a = o4_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_135 =>
            -- reg_a = o5_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_136 =>
            -- reg_a = a0_X; reg_b = a7_X; reg_acc = reg_o; o7_X = reg_o; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "111";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_137 =>
            -- reg_a = a1_X; reg_b = a7_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_138 =>
            -- reg_a = o1_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_139 =>
            -- reg_a = a2_X; reg_b = a6_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_140 =>
            -- reg_a = o2_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_141 =>
            -- reg_a = a3_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_142 =>
            -- reg_a = o3_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_143 =>
            -- reg_a = a4_X; reg_b = a4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_144 =>
            -- reg_a = o4_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_145 =>
            -- reg_a = o5_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_146 =>
            -- reg_a = o6_X; reg_b = primeSP2; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_147 =>
            -- reg_a = a2_X; reg_b = a7_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_148 =>
            -- reg_a = o2_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_149 =>
            -- reg_a = a3_X; reg_b = a6_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_150 =>
            -- reg_a = o3_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_151 =>
            -- reg_a = a4_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_152 =>
            -- reg_a = o4_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_153 =>
            -- reg_a = o5_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_154 =>
            -- reg_a = o6_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_155 =>
            -- reg_a = o7_X; reg_b = primeSP2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_156 =>
            -- reg_a = a3_X; reg_b = a7_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_157 =>
            -- reg_a = o3_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_158 =>
            -- reg_a = a4_X; reg_b = a6_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_159 =>
            -- reg_a = o4_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_160 =>
            -- reg_a = a5_X; reg_b = a5_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_161 =>
            -- reg_a = o5_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_162 =>
            -- reg_a = o6_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_163 =>
            -- reg_a = o7_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_164 =>
            -- reg_a = a4_X; reg_b = a7_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_165 =>
            -- reg_a = o4_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_166 =>
            -- reg_a = a5_X; reg_b = a6_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_167 =>
            -- reg_a = o5_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_168 =>
            -- reg_a = o6_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_169 =>
            -- reg_a = o7_X; reg_b = primeSP4; reg_acc = reg_o; o3_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_170 =>
            -- reg_a = a5_X; reg_b = a7_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_171 =>
            -- reg_a = o5_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_172 =>
            -- reg_a = a6_X; reg_b = a6_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_173 =>
            -- reg_a = o6_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_174 =>
            -- reg_a = o7_X; reg_b = primeSP5; reg_acc = reg_o; o4_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_175 =>
            -- reg_a = a6_X; reg_b = a7_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_176 =>
            -- reg_a = o6_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_177 =>
            -- reg_a = o7_X; reg_b = primeSP6; reg_acc = reg_o; o5_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_178 =>
            -- reg_a = a7_X; reg_b = a7_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_179 =>
            -- reg_a = o7_X; reg_b = primeSP7; reg_acc = reg_o; o6_X = reg_o; o7_X = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_0 =>
            -- -- In case of sizes 3, 4, 5, 6, 7, 8
            -- reg_a = a0_X; reg_b = a0_X; reg_acc = 0; o0_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_1 =>
            -- reg_a = a0_X; reg_b = a1_X; reg_acc = reg_o >> 256; o1_X = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_2 =>
            -- reg_a = a1_X; reg_b = a1_X; reg_acc = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_3 =>
            -- -- In case of size 3
            -- reg_a = a0_X; reg_b = a2_X; reg_acc = reg_o; o2_X = reg_o; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_4 =>
            -- reg_a = a1_X; reg_b = a2_X; reg_acc = reg_o >> 256; Enable sign b; o0_X = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_5 =>
            -- reg_a = a2_X; reg_b = a2_X; reg_acc = reg_o >> 256; Enable sign a,b; o1_X = reg_o; o2_X = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_7 =>
            -- -- In case of sizes 4, 5, 6, 7, 8
            -- reg_a = a0_X; reg_b = a2_X; reg_acc = reg_o; o2_X = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_8 =>
            -- reg_a = o0_X; reg_b = primeSP3; reg_acc = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_9 =>
            -- reg_a = a1_X; reg_b = a2_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_10 =>
            -- -- In case of size 4
            -- reg_a = a0_X; reg_b = a3_X; reg_acc = reg_o; o3_X = reg_o; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_11 =>
            -- reg_a = a1_X; reg_b = a3_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_12 =>
            -- reg_a = o1_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_13 =>
            -- reg_a = a2_X; reg_b = a2_X; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_14 =>
            -- reg_a = a2_X; reg_b = a3_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_15 =>
            -- reg_a = o2_X; reg_b = primeSP3; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_16 =>
            -- reg_a = a3_X; reg_b = a3_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_17 =>
            -- reg_a = o3_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; o3_X = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_19 =>
            -- -- In case of sizes 5, 6, 7, 8
            -- reg_a = a0_X; reg_b = a3_X; reg_acc = reg_o; o3_X = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_20 =>
            -- reg_a = o0_X; reg_b = primeSP4; reg_acc = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_21 =>
            -- reg_a = a1_X; reg_b = a3_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_22 =>
            -- reg_a = o1_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_23 =>
            -- reg_a = a2_X; reg_b = a2_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_24 =>
            -- -- In case of size 5
            -- reg_a = a0_X; reg_b = a4_X; reg_acc = reg_o; o4_X = reg_o; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_25 =>
            -- reg_a = a1_X; reg_b = a4_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_26 =>
            -- reg_a = o1_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_27 =>
            -- reg_a = a2_X; reg_b = a3_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_28 =>
            -- reg_a = o2_X; reg_b = primeSP3; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_29 =>
            -- reg_a = a2_X; reg_b = a4_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_30 =>
            -- reg_a = o2_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_31 =>
            -- reg_a = a3_X; reg_b = a3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_32 =>
            -- reg_a = o3_X; reg_b = primeSP3; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_33 =>
            -- reg_a = a3_X; reg_b = a4_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_34 =>
            -- reg_a = o3_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_35 =>
            -- reg_a = o4_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_36 =>
            -- reg_a = a4_X; reg_b = a4_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_37 =>
            -- reg_a = o4_X; reg_b = primeSP4; reg_acc = reg_o; o3_X = reg_o; o4_X = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_39 =>
            -- -- In case of sizes 6, 7, 8
            -- reg_a = a0_X; reg_b = a4_X; reg_acc = reg_o; o4_X = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_40 =>
            -- reg_a = o0_X; reg_b = primeSP5; reg_acc = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_41 =>
            -- reg_a = a1_X; reg_b = a4_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_42 =>
            -- reg_a = o1_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_43 =>
            -- reg_a = a2_X; reg_b = a3_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_44 =>
            -- reg_a = o2_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_45 =>
            -- -- In case of size 6
            -- reg_a = a0_X; reg_b = a5_X; reg_acc = reg_o; o5_X = reg_o; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_46 =>
            -- reg_a = a1_X; reg_b = a5_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_47 =>
            -- reg_a = o1_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_48 =>
            -- reg_a = a2_X; reg_b = a4_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_49 =>
            -- reg_a = o2_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_50 =>
            -- reg_a = a3_X; reg_b = a3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_51 =>
            -- reg_a = o3_X; reg_b = primeSP3; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_52 =>
            -- reg_a = a2_X; reg_b = a5_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_53 =>
            -- reg_a = o2_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_54 =>
            -- reg_a = a3_X; reg_b = a4_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_55 =>
            -- reg_a = o3_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_56 =>
            -- reg_a = o4_X; reg_b = primeSP3; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_57 =>
            -- reg_a = a3_X; reg_b = a5_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_58 =>
            -- reg_a = o3_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_59 =>
            -- reg_a = a4_X; reg_b = a4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_60 =>
            -- reg_a = o4_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_61 =>
            -- reg_a = o5_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_62 =>
            -- reg_a = a4_X; reg_b = a5_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_63 =>
            -- reg_a = o4_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_64 =>
            -- reg_a = o5_X; reg_b = primeSP4; reg_acc = reg_o; o3_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_65 =>
            -- reg_a = a5_X; reg_b = a5_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_66 =>
            -- reg_a = o5_X; reg_b = primeSP5; reg_acc = reg_o; o4_X = reg_o; o5_X = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_68 =>
            -- -- In case of sizes 7, 8
            -- reg_a = a0_X; reg_b = a5_X; reg_acc = reg_o; o5_X = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_69 =>
            -- reg_a = o0_X; reg_b = primeSP6; reg_acc = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_70 =>
            -- reg_a = a1_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_71 =>
            -- reg_a = o1_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_72 =>
            -- reg_a = a2_X; reg_b = a4_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_73 =>
            -- reg_a = o2_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_74 =>
            -- reg_a = a3_X; reg_b = a3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_75 =>
            -- reg_a = o3_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_76 =>
            -- -- In case of size 7
            -- reg_a = a0_X; reg_b = a6_X; reg_acc = reg_o; o6_X = reg_o; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_77 =>
            -- reg_a = a1_X; reg_b = a6_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_78 =>
            -- reg_a = o1_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_79 =>
            -- reg_a = a2_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_80 =>
            -- reg_a = o2_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_81 =>
            -- reg_a = a3_X; reg_b = a4_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_82 =>
            -- reg_a = o3_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_83 =>
            -- reg_a = o4_X; reg_b = primeSP3; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_84 =>
            -- reg_a = a2_X; reg_b = a6_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_85 =>
            -- reg_a = o2_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_86 =>
            -- reg_a = a3_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_87 =>
            -- reg_a = o3_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_88 =>
            -- reg_a = a4_X; reg_b = a4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_89 =>
            -- reg_a = o4_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_90 =>
            -- reg_a = o5_X; reg_b = primeSP3; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_91 =>
            -- reg_a = a3_X; reg_b = a6_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_92 =>
            -- reg_a = o3_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_93 =>
            -- reg_a = a4_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_94 =>
            -- reg_a = o4_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_95 =>
            -- reg_a = o5_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_96 =>
            -- reg_a = o6_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_97 =>
            -- reg_a = a4_X; reg_b = a6_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_98 =>
            -- reg_a = o4_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_99 =>
            -- reg_a = a5_X; reg_b = a5_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_100 =>
            -- reg_a = o5_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_101 =>
            -- reg_a = o6_X; reg_b = primeSP4; reg_acc = reg_o; o3_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_102 =>
            -- reg_a = a5_X; reg_b = a6_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_103 =>
            -- reg_a = o5_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_104 =>
            -- reg_a = o6_X; reg_b = primeSP5; reg_acc = reg_o; o4_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_105 =>
            -- reg_a = a6_X; reg_b = a6_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_106 =>
            -- reg_a = o6_X; reg_b = primeSP6; reg_acc = reg_o; o5_X = reg_o; o6_X = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_108 =>
            -- -- In case of size 8
            -- reg_a = a0_X; reg_b = a6_X; reg_acc = reg_o; o6_X = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_109 =>
            -- reg_a = o0_X; reg_b = primeSP7; reg_acc = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_110 =>
            -- reg_a = a1_X; reg_b = a6_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_111 =>
            -- reg_a = o1_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_112 =>
            -- reg_a = a2_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_113 =>
            -- reg_a = o2_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_114 =>
            -- reg_a = a3_X; reg_b = a4_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_115 =>
            -- reg_a = o3_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_116 =>
            -- reg_a = o4_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_117 =>
            -- reg_a = a0_X; reg_b = a7_X; reg_acc = reg_o; o7_X = reg_o; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "111";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_118 =>
            -- reg_a = a1_X; reg_b = a7_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_119 =>
            -- reg_a = o1_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_120 =>
            -- reg_a = a2_X; reg_b = a6_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_121 =>
            -- reg_a = o2_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_122 =>
            -- reg_a = a3_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_123 =>
            -- reg_a = o3_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_124 =>
            -- reg_a = a4_X; reg_b = a4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_125 =>
            -- reg_a = o4_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_126 =>
            -- reg_a = o5_X; reg_b = primeSP3; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_127 =>
            -- reg_a = a2_X; reg_b = a7_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_128 =>
            -- reg_a = o2_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_129 =>
            -- reg_a = a3_X; reg_b = a6_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_130 =>
            -- reg_a = o3_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_131 =>
            -- reg_a = a4_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_132 =>
            -- reg_a = o4_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_133 =>
            -- reg_a = o5_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_134 =>
            -- reg_a = o6_X; reg_b = primeSP3; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_135 =>
            -- reg_a = a3_X; reg_b = a7_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_136 =>
            -- reg_a = o3_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_137 =>
            -- reg_a = a4_X; reg_b = a6_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_138 =>
            -- reg_a = o4_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_139 =>
            -- reg_a = a5_X; reg_b = a5_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_140 =>
            -- reg_a = o5_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_141 =>
            -- reg_a = o6_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_142 =>
            -- reg_a = o7_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_143 =>
            -- reg_a = a4_X; reg_b = a7_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_144 =>
            -- reg_a = o4_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_145 =>
            -- reg_a = a5_X; reg_b = a6_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_146 =>
            -- reg_a = o5_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_147 =>
            -- reg_a = o6_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_148 =>
            -- reg_a = o7_X; reg_b = primeSP4; reg_acc = reg_o; o3_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_149 =>
            -- reg_a = a5_X; reg_b = a7_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_150 =>
            -- reg_a = o5_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_151 =>
            -- reg_a = a6_X; reg_b = a6_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_152 =>
            -- reg_a = o6_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_153 =>
            -- reg_a = o7_X; reg_b = primeSP5; reg_acc = reg_o; o4_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_154 =>
            -- reg_a = a6_X; reg_b = a7_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_155 =>
            -- reg_a = o6_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_156 =>
            -- reg_a = o7_X; reg_b = primeSP6; reg_acc = reg_o; o5_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_157 =>
            -- reg_a = a7_X; reg_b = a7_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_158 =>
            -- reg_a = o7_X; reg_b = primeSP7; reg_acc = reg_o; o6_X = reg_o; o7_X = reg_o >> 256; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_direct_0 =>
            -- -- In case of size 1
            -- reg_a = a0_X; reg_b = b0_X; reg_acc = 0; o0_0 = reg_o; Enable sign a,b; operation : b +/- a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '1';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_direct_2 =>
            -- -- In case of size 2, 3, 4, 5, 6, 7, 8
            -- reg_a = a0_X; reg_b = b0_X; reg_acc = 0; o0_X = reg_o; operation : b +/- a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '1';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_direct_3 =>
            -- -- In case of size 2
            -- reg_a = a1_X; reg_b = b1_X; reg_acc = reg_o >> 256; o1_X = reg_o; Enable sign a, b; operation : b +/- a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '1';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_direct_5 =>
            -- -- In case of size 3, 4, 5, 6, 7, 8
            -- reg_a = a1_X; reg_b = b1_X; reg_acc = reg_o >> 256; o1_X = reg_o; operation : b +/- a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '1';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_direct_6 =>
            -- -- In case of size 3
            -- reg_a = a2_X; reg_b = b2_X; reg_acc = reg_o >> 256; o2_X = reg_o; Enable sign a,b; operation : b +/- a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '1';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_direct_8 =>
            -- -- In case of size 4, 5, 6, 7, 8
            -- reg_a = a2_X; reg_b = b2_X; reg_acc = reg_o >> 256; o2_X = reg_o; operation : b +/- a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '1';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_direct_9 =>
            -- -- In case of size 4
            -- reg_a = a3_X; reg_b = b3_X; reg_acc = reg_o >> 256; o3_X = reg_o; Enable sign a,b; operation : b +/- a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '1';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_direct_11 =>
            -- -- In case of size 4, 5, 6, 7, 8
            -- reg_a = a3_X; reg_b = b3_X; reg_acc = reg_o >> 256; o3_X = reg_o; operation : b +/- a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '1';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_direct_12 =>
            -- -- In case of size 5
            -- reg_a = a4_X; reg_b = b4_X; reg_acc = reg_o >> 256; o4_X = reg_o; Enable sign a,b; operation : b +/- a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '1';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_direct_14 =>
            -- -- In case of size 6, 7, 8
            -- reg_a = a4_X; reg_b = b4_X; reg_acc = reg_o >> 256; o4_X = reg_o; operation : b +/- a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '1';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_direct_15 =>
            -- -- In case of size 6
            -- reg_a = a5_X; reg_b = b5_X; reg_acc = reg_o >> 256; o5_X = reg_o; Enable sign a,b; operation : b +/- a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '1';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_direct_17 =>
            -- -- In case of size 7, 8
            -- reg_a = a5_X; reg_b = b5_X; reg_acc = reg_o >> 256; o5_X = reg_o; operation : b +/- a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '1';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_direct_18 =>
            -- -- In case of size 7
            -- reg_a = a6_X; reg_b = b6_X; reg_acc = reg_o >> 256; o6_X = reg_o; Enable sign a,b; operation : b +/- a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '1';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_direct_20 =>
            -- -- In case of size 8
            -- reg_a = a6_X; reg_b = b6_X; reg_acc = reg_o >> 256; o6_X = reg_o; operation : b +/- a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '1';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_direct_21 =>
            -- reg_a = a7_X; reg_b = b7_X; reg_acc = reg_o >> 256; o7_X = reg_o; Enable sign a,b; operation : b +/- a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "111";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '1';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_0 =>
            -- -- In case of size 1
            -- reg_a = a0_X; reg_b = 0; reg_acc = 0; Enable sign a,b; operation : b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '1';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_1 =>
            -- reg_a = 0; reg_b = prime0; reg_acc = reg_o; reg_s = reg_o_positive; Enable sign a,b; operation : -s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "11";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '1';
            next_mac_sel_reg_s_reg_o_sign <= '1';
            next_mac_reg_s_reg_o_positive <= '1';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_2 =>
            -- reg_a = 0; reg_b = prime0; reg_acc = reg_o; reg_s = reg_o_negative; Enable sign a,b; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "11";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '1';
            next_mac_sel_reg_s_reg_o_sign <= '1';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_3 =>
            -- reg_a = 0; reg_b = prime0; reg_acc = reg_o; o0_X = reg_o; reg_s = reg_o_negative; Enable sign a,b; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "11";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '1';
            next_mac_sel_reg_s_reg_o_sign <= '1';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_5 =>
            -- -- In case of size 2
            -- reg_a = a1_X; reg_b = 0; reg_acc = 0; Enable sign a,b; operation : b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '1';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_6 =>
            -- reg_a = a0_X; reg_b = prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_positive; operation : -s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '1';
            next_mac_sel_reg_s_reg_o_sign <= '1';
            next_mac_reg_s_reg_o_positive <= '1';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_7 =>
            -- reg_a = a1_X; reg_b = prime1; reg_acc = reg_o >> 256; o1_X = reg_o; Enable sign a,b; operation : -s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_8 =>
            -- reg_a = o0_X; reg_b = prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '1';
            next_mac_sel_reg_s_reg_o_sign <= '1';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_9 =>
            -- reg_a = o1_X; reg_b = prime1; reg_acc = reg_o >> 256; o1_X = reg_o; Enable sign a,b operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_10 =>
            -- reg_a = o0_X; reg_b = prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '1';
            next_mac_sel_reg_s_reg_o_sign <= '1';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_11 =>
            -- reg_a = o1_X; reg_b = prime1; reg_acc = reg_o >> 256; o1_X = reg_o; Enable sign a,b operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_13 =>
            -- -- In case of size 3
            -- reg_a = a2_X; reg_b = 0; reg_acc = 0; Enable sign a,b; operation : b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '1';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_14 =>
            -- reg_a = a0_X; reg_b = prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_positive; operation : -s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '1';
            next_mac_sel_reg_s_reg_o_sign <= '1';
            next_mac_reg_s_reg_o_positive <= '1';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_15 =>
            -- reg_a = a1_X; reg_b = prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : -s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_16 =>
            -- reg_a = a2_X; reg_b = prime2; reg_acc = reg_o >> 256; o2_X = reg_o; Enable sign a,b; operation : -s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_17 =>
            -- reg_a = o0_X; reg_b = prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '1';
            next_mac_sel_reg_s_reg_o_sign <= '1';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_18 =>
            -- reg_a = o1_X; reg_b = prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_19 =>
            -- reg_a = o2_X; reg_b = prime2; reg_acc = reg_o >> 256; o2_X = reg_o; Enable sign a,b operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_20 =>
            -- reg_a = o0_X; reg_b = prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '1';
            next_mac_sel_reg_s_reg_o_sign <= '1';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_21 =>
            -- reg_a = o1_X; reg_b = prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_22 =>
            -- reg_a = o2_X; reg_b = prime2; reg_acc = reg_o >> 256; o2_X = reg_o; Enable sign a,b operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_24 =>
            -- -- In case of size 4
            -- reg_a = a3_X; reg_b = 0; reg_acc = 0; Enable sign a,b; operation : b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '1';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_25 =>
            -- reg_a = a0_X; reg_b = prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_positive; operation : -s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '1';
            next_mac_sel_reg_s_reg_o_sign <= '1';
            next_mac_reg_s_reg_o_positive <= '1';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_26 =>
            -- reg_a = a1_X; reg_b = prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : -s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_27 =>
            -- reg_a = a2_X; reg_b = prime2; reg_acc = reg_o >> 256; o2_X = reg_o; operation : -s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_28 =>
            -- reg_a = a3_X; reg_b = prime3; reg_acc = reg_o >> 256; o3_X = reg_o; Enable sign a,b; operation : -s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_29 =>
            -- reg_a = o0_X; reg_b = prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '1';
            next_mac_sel_reg_s_reg_o_sign <= '1';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_30 =>
            -- reg_a = o1_X; reg_b = prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_31 =>
            -- reg_a = o2_X; reg_b = prime2; reg_acc = reg_o >> 256; o2_X = reg_o; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_32 =>
            -- reg_a = o3_X; reg_b = prime3; reg_acc = reg_o >> 256; o3_X = reg_o; Enable sign a,b; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_33 =>
            -- reg_a = o0_X; reg_b = prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '1';
            next_mac_sel_reg_s_reg_o_sign <= '1';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_34 =>
            -- reg_a = o1_X; reg_b = prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_35 =>
            -- reg_a = o2_X; reg_b = prime2; reg_acc = reg_o >> 256; o2_X = reg_o; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_36 =>
            -- reg_a = o3_X; reg_b = prime3; reg_acc = reg_o >> 256; o3_X = reg_o; Enable sign a,b; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_38 =>
            -- -- In case of size 5
            -- reg_a = a4_X; reg_b = 0; reg_acc = 0; Enable sign a,b; operation : b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '1';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_39 =>
            -- reg_a = a0_X; reg_b = prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_positive; operation : -s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '1';
            next_mac_sel_reg_s_reg_o_sign <= '1';
            next_mac_reg_s_reg_o_positive <= '1';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_40 =>
            -- reg_a = a1_X; reg_b = prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : -s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_41 =>
            -- reg_a = a2_X; reg_b = prime2; reg_acc = reg_o >> 256; o2_X = reg_o; operation : -s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_42 =>
            -- reg_a = a3_X; reg_b = prime3; reg_acc = reg_o >> 256; o3_X = reg_o; operation : -s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_43 =>
            -- reg_a = a4_X; reg_b = prime4; reg_acc = reg_o >> 256; o4_X = reg_o; Enable sign a,b; operation : -s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_44 =>
            -- reg_a = o0_X; reg_b = prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '1';
            next_mac_sel_reg_s_reg_o_sign <= '1';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_45 =>
            -- reg_a = o1_X; reg_b = prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_46 =>
            -- reg_a = o2_X; reg_b = prime2; reg_acc = reg_o >> 256; o2_X = reg_o; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_47 =>
            -- reg_a = o3_X; reg_b = prime3; reg_acc = reg_o >> 256; o3_X = reg_o; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_48 =>
            -- reg_a = o4_X; reg_b = prime4; reg_acc = reg_o >> 256; o4_X = reg_o; Enable sign a,b; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_49 =>
            -- reg_a = o0_X; reg_b = prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '1';
            next_mac_sel_reg_s_reg_o_sign <= '1';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_50 =>
            -- reg_a = o1_X; reg_b = prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_51 =>
            -- reg_a = o2_X; reg_b = prime2; reg_acc = reg_o >> 256; o2_X = reg_o; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_52 =>
            -- reg_a = o3_X; reg_b = prime3; reg_acc = reg_o >> 256; o3_X = reg_o; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_53 =>
            -- reg_a = o4_X; reg_b = prime4; reg_acc = reg_o >> 256; o4_X = reg_o; Enable sign a,b; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_55 =>
            -- -- In case of size 6
            -- reg_a = a5_X; reg_b = 0; reg_acc = 0; Enable sign a,b; operation : b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '1';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_56 =>
            -- reg_a = a0_X; reg_b = prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_positive; operation : -s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '1';
            next_mac_sel_reg_s_reg_o_sign <= '1';
            next_mac_reg_s_reg_o_positive <= '1';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_57 =>
            -- reg_a = a1_X; reg_b = prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : -s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_58 =>
            -- reg_a = a2_X; reg_b = prime2; reg_acc = reg_o >> 256; o2_X = reg_o; operation : -s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_59 =>
            -- reg_a = a3_X; reg_b = prime3; reg_acc = reg_o >> 256; o3_X = reg_o; operation : -s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_60 =>
            -- reg_a = a4_X; reg_b = prime4; reg_acc = reg_o >> 256; o4_X = reg_o; operation : -s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_61 =>
            -- reg_a = a5_X; reg_b = prime5; reg_acc = reg_o >> 256; o5_X = reg_o; Enable sign a,b; operation : -s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_62 =>
            -- reg_a = o0_X; reg_b = prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '1';
            next_mac_sel_reg_s_reg_o_sign <= '1';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_63 =>
            -- reg_a = o1_X; reg_b = prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_64 =>
            -- reg_a = o2_X; reg_b = prime2; reg_acc = reg_o >> 256; o2_X = reg_o; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_65 =>
            -- reg_a = o3_X; reg_b = prime3; reg_acc = reg_o >> 256; o3_X = reg_o; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_66 =>
            -- reg_a = o4_X; reg_b = prime4; reg_acc = reg_o >> 256; o4_X = reg_o; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_67 =>
            -- reg_a = o5_X; reg_b = prime5; reg_acc = reg_o >> 256; o5_X = reg_o; Enable sign a,b; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_68 =>
            -- reg_a = o0_X; reg_b = prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '1';
            next_mac_sel_reg_s_reg_o_sign <= '1';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_69 =>
            -- reg_a = o1_X; reg_b = prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_70 =>
            -- reg_a = o2_X; reg_b = prime2; reg_acc = reg_o >> 256; o2_X = reg_o; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_71 =>
            -- reg_a = o3_X; reg_b = prime3; reg_acc = reg_o >> 256; o3_X = reg_o; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_72 =>
            -- reg_a = o4_X; reg_b = prime4; reg_acc = reg_o >> 256; o4_X = reg_o; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_73 =>
            -- reg_a = o5_X; reg_b = prime5; reg_acc = reg_o >> 256; o5_X = reg_o; Enable sign a,b; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_75 =>
            -- -- In case of size 7
            -- reg_a = a6_X; reg_b = 0; reg_acc = 0; Enable sign a,b; operation : b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '1';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_76 =>
            -- reg_a = a0_X; reg_b = prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_positive; operation : -s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '1';
            next_mac_sel_reg_s_reg_o_sign <= '1';
            next_mac_reg_s_reg_o_positive <= '1';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_77 =>
            -- reg_a = a1_X; reg_b = prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : -s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_78 =>
            -- reg_a = a2_X; reg_b = prime2; reg_acc = reg_o >> 256; o2_X = reg_o; operation : -s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_79 =>
            -- reg_a = a3_X; reg_b = prime3; reg_acc = reg_o >> 256; o3_X = reg_o; operation : -s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_80 =>
            -- reg_a = a4_X; reg_b = prime4; reg_acc = reg_o >> 256; o4_X = reg_o; operation : -s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_81 =>
            -- reg_a = a5_X; reg_b = prime5; reg_acc = reg_o >> 256; o5_X = reg_o; operation : -s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_82 =>
            -- reg_a = a6_X; reg_b = prime6; reg_acc = reg_o >> 256; o6_X = reg_o; Enable sign a,b; operation : -s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_83 =>
            -- reg_a = o0_X; reg_b = prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '1';
            next_mac_sel_reg_s_reg_o_sign <= '1';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_84 =>
            -- reg_a = o1_X; reg_b = prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_85 =>
            -- reg_a = o2_X; reg_b = prime2; reg_acc = reg_o >> 256; o2_X = reg_o; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_86 =>
            -- reg_a = o3_X; reg_b = prime3; reg_acc = reg_o >> 256; o3_X = reg_o; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_87 =>
            -- reg_a = o4_X; reg_b = prime4; reg_acc = reg_o >> 256; o4_X = reg_o; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_88 =>
            -- reg_a = o5_X; reg_b = prime5; reg_acc = reg_o >> 256; o5_X = reg_o; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_89 =>
            -- reg_a = o6_X; reg_b = prime6; reg_acc = reg_o >> 256; o6_X = reg_o; Enable sign a,b; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_90 =>
            -- reg_a = o0_X; reg_b = prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '1';
            next_mac_sel_reg_s_reg_o_sign <= '1';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_91 =>
            -- reg_a = o1_X; reg_b = prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_92 =>
            -- reg_a = o2_X; reg_b = prime2; reg_acc = reg_o >> 256; o2_X = reg_o; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_93 =>
            -- reg_a = o3_X; reg_b = prime3; reg_acc = reg_o >> 256; o3_X = reg_o; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_94 =>
            -- reg_a = o4_X; reg_b = prime4; reg_acc = reg_o >> 256; o4_X = reg_o; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_95 =>
            -- reg_a = o5_X; reg_b = prime5; reg_acc = reg_o >> 256; o5_X = reg_o; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_96 =>
            -- reg_a = o6_X; reg_b = prime6; reg_acc = reg_o >> 256; o6_X = reg_o; Enable sign a,b; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_98 =>
            -- -- In case of size 8
            -- reg_a = a7_X; reg_b = 0; reg_acc = 0; Enable sign a,b; operation : b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "111";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '1';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_99 =>
            -- reg_a = a0_X; reg_b = prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_positive; operation : -s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '1';
            next_mac_sel_reg_s_reg_o_sign <= '1';
            next_mac_reg_s_reg_o_positive <= '1';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_100 =>
            -- reg_a = a1_X; reg_b = prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : -s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_101 =>
            -- reg_a = a2_X; reg_b = prime2; reg_acc = reg_o >> 256; o2_X = reg_o; operation : -s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_102 =>
            -- reg_a = a3_X; reg_b = prime3; reg_acc = reg_o >> 256; o3_X = reg_o; operation : -s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_103 =>
            -- reg_a = a4_X; reg_b = prime4; reg_acc = reg_o >> 256; o4_X = reg_o; operation : -s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_104 =>
            -- reg_a = a5_X; reg_b = prime5; reg_acc = reg_o >> 256; o5_X = reg_o; operation : -s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_105 =>
            -- reg_a = a6_X; reg_b = prime6; reg_acc = reg_o >> 256; o6_X = reg_o; operation : -s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_106 =>
            -- reg_a = a7_X; reg_b = prime7; reg_acc = reg_o >> 256; o7_X = reg_o; Enable sign a,b; operation : -s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "111";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_107 =>
            -- reg_a = o0_X; reg_b = prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '1';
            next_mac_sel_reg_s_reg_o_sign <= '1';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_108 =>
            -- reg_a = o1_X; reg_b = prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_109 =>
            -- reg_a = o2_X; reg_b = prime2; reg_acc = reg_o >> 256; o2_X = reg_o; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_110 =>
            -- reg_a = o3_X; reg_b = prime3; reg_acc = reg_o >> 256; o3_X = reg_o; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_111 =>
            -- reg_a = o4_X; reg_b = prime4; reg_acc = reg_o >> 256; o4_X = reg_o; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_112 =>
            -- reg_a = o5_X; reg_b = prime5; reg_acc = reg_o >> 256; o5_X = reg_o; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_113 =>
            -- reg_a = o6_X; reg_b = prime6; reg_acc = reg_o >> 256; o6_X = reg_o; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_114 =>
            -- reg_a = o7_X; reg_b = prime7; reg_acc = reg_o >> 256; o7_X = reg_o; Enable sign a,b; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "111";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_115 =>
            -- reg_a = o0_X; reg_b = prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '1';
            next_mac_sel_reg_s_reg_o_sign <= '1';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_116 =>
            -- reg_a = o1_X; reg_b = prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_117 =>
            -- reg_a = o2_X; reg_b = prime2; reg_acc = reg_o >> 256; o2_X = reg_o; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_118 =>
            -- reg_a = o3_X; reg_b = prime3; reg_acc = reg_o >> 256; o3_X = reg_o; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_119 =>
            -- reg_a = o4_X; reg_b = prime4; reg_acc = reg_o >> 256; o4_X = reg_o; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_120 =>
            -- reg_a = o5_X; reg_b = prime5; reg_acc = reg_o >> 256; o5_X = reg_o; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_121 =>
            -- reg_a = o6_X; reg_b = prime6; reg_acc = reg_o >> 256; o6_X = reg_o; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_122 =>
            -- reg_a = o7_X; reg_b = prime7; reg_acc = reg_o >> 256; o7_X = reg_o; Enable sign a,b; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "111";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_0 =>
            -- Operands size 1
            -- reg_a = a0_X; reg_b = b0_X; reg_acc = 0; o0_X = reg_o; Enable sign a,b; operation : b +/- a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '1';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_1 =>
            -- reg_a = 0; reg_b = 2prime0; reg_acc = reg_o; reg_s = reg_o_positive; o0_X = reg_o; Enable sign a,b; operation : -s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "11";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '1';
            next_mac_sel_reg_s_reg_o_sign <= '1';
            next_mac_reg_s_reg_o_positive <= '1';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_2 =>
            -- reg_a = 0; reg_b = 2prime0; reg_acc = reg_o; reg_s = reg_o_negative; o0_X = reg_o; Enable sign a,b; operation : s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "11";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '1';
            next_mac_sel_reg_s_reg_o_sign <= '1';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_3 =>
            -- reg_a = 0; reg_b = 2prime0; reg_acc = reg_o; reg_s = reg_o_negative; o0_X = reg_o; Enable sign a,b; operation : s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "11";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '1';
            next_mac_sel_reg_s_reg_o_sign <= '1';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_5 =>
            -- -- In case of sizes 2, 3, 4, 5, 6, 7, 8
            -- reg_a = a0_X; reg_b = b0_X; reg_acc = 0; o0_X = reg_o; operation : b +/- a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '1';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_6 =>
            -- -- In case of size 2
            -- reg_a = a1_X; reg_b = b1_X; reg_acc = reg_o >> 256; o1_X = reg_o; Enable sign a, b; operation : b +/- a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '1';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_7 =>
            -- reg_a = o0_X; reg_b = 2prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_positive; operation : -s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '1';
            next_mac_sel_reg_s_reg_o_sign <= '1';
            next_mac_reg_s_reg_o_positive <= '1';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_8 =>
            -- reg_a = o1_X; reg_b = 2prime1; reg_acc = reg_o >> 256; o1_X = reg_o; Enable sign a,b; operation : -s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_9 =>
            -- reg_a = o0_X; reg_b = 2prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '1';
            next_mac_sel_reg_s_reg_o_sign <= '1';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_10 =>
            -- reg_a = o1_X; reg_b = 2prime1; reg_acc = reg_o >> 256; o1_X = reg_o; Enable sign a,b; operation : s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_11 =>
            -- reg_a = o0_X; reg_b = 2prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '1';
            next_mac_sel_reg_s_reg_o_sign <= '1';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_12 =>
            -- reg_a = o1_X; reg_b = 2prime1; reg_acc = reg_o >> 256; o1_X = reg_o; Enable sign a,b; operation : s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_14 =>
            -- -- In case of sizes 3, 4, 5, 6, 7, 8
            -- reg_a = a1_X; reg_b = b1_X; reg_acc = reg_o >> 256; o1_X = reg_o; operation : b +/- a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '1';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_15 =>
            -- -- In case of size 3
            -- reg_a = a2_X; reg_b = b2_X; reg_acc = reg_o >> 256; o2_X = reg_o; Enable sign a, b; operation : b +/- a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '1';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_16 =>
            -- reg_a = o0_X; reg_b = 2prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_positive; operation : -s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '1';
            next_mac_sel_reg_s_reg_o_sign <= '1';
            next_mac_reg_s_reg_o_positive <= '1';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_17 =>
            -- reg_a = o1_X; reg_b = 2prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : -s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_18 =>
            -- reg_a = o2_X; reg_b = 2prime2; reg_acc = reg_o >> 256; o2_X = reg_o; Enable sign a,b; operation : -s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_19 =>
            -- reg_a = o0_X; reg_b = 2prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '1';
            next_mac_sel_reg_s_reg_o_sign <= '1';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_20 =>
            -- reg_a = o1_X; reg_b = 2prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_21 =>
            -- reg_a = o2_X; reg_b = 2prime2; reg_acc = reg_o >> 256; o2_X = reg_o; Enable sign a,b; operation : s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_22 =>
            -- reg_a = o0_X; reg_b = 2prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '1';
            next_mac_sel_reg_s_reg_o_sign <= '1';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_23 =>
            -- reg_a = o1_X; reg_b = 2prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_24 =>
            -- reg_a = o2_X; reg_b = 2prime2; reg_acc = reg_o >> 256; o2_X = reg_o; Enable sign a,b; operation : s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_26 =>
            -- -- In case of size 4, 5, 6, 7, 8
            -- reg_a = a2_X; reg_b = b2_X; reg_acc = reg_o >> 256; o2_X = reg_o; operation : b +/- a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '1';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_27 =>
            -- -- In case of size 4
            -- reg_a = a3_X; reg_b = b3_X; reg_acc = reg_o >> 256; o3_X = reg_o; Enable sign a, b; operation : b +/- a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '1';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_28 =>
            -- reg_a = o0_X; reg_b = 2prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_positive; operation : -s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '1';
            next_mac_sel_reg_s_reg_o_sign <= '1';
            next_mac_reg_s_reg_o_positive <= '1';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_29 =>
            -- reg_a = o1_X; reg_b = 2prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : -s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_30 =>
            -- reg_a = o2_X; reg_b = 2prime2; reg_acc = reg_o >> 256; o2_X = reg_o; operation : -s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_31 =>
            -- reg_a = o3_X; reg_b = 2prime3; reg_acc = reg_o >> 256; o3_X = reg_o; Enable sign a,b; operation : -s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_32 =>
            -- reg_a = o0_X; reg_b = 2prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '1';
            next_mac_sel_reg_s_reg_o_sign <= '1';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_33 =>
            -- reg_a = o1_X; reg_b = 2prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_34 =>
            -- reg_a = o2_X; reg_b = 2prime2; reg_acc = reg_o >> 256; o2_X = reg_o; operation : s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_35 =>
            -- reg_a = o3_X; reg_b = 2prime3; reg_acc = reg_o >> 256; o3_X = reg_o; Enable sign a,b; operation : s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_36 =>
            -- reg_a = o0_X; reg_b = 2prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '1';
            next_mac_sel_reg_s_reg_o_sign <= '1';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_37 =>
            -- reg_a = o1_X; reg_b = 2prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_38 =>
            -- reg_a = o2_X; reg_b = 2prime2; reg_acc = reg_o >> 256; o2_X = reg_o; operation : s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_39 =>
            -- reg_a = o3_X; reg_b = 2prime3; reg_acc = reg_o >> 256; o3_X = reg_o; Enable sign a,b; operation : s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_41 =>
            -- -- In case of size 5, 6, 7, 8
            -- reg_a = a3_X; reg_b = b3_X; reg_acc = reg_o >> 256; o3_X = reg_o; operation : b +/- a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '1';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_42 =>
            -- -- In case of size 5
            -- reg_a = a4_X; reg_b = b4_X; reg_acc = reg_o >> 256; o4_X = reg_o; Enable sign a, b; operation : b +/- a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '1';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_43 =>
            -- reg_a = o0_X; reg_b = 2prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_positive; operation : -s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '1';
            next_mac_sel_reg_s_reg_o_sign <= '1';
            next_mac_reg_s_reg_o_positive <= '1';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_44 =>
            -- reg_a = o1_X; reg_b = 2prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : -s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_45 =>
            -- reg_a = o2_X; reg_b = 2prime2; reg_acc = reg_o >> 256; o2_X = reg_o; operation : -s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_46 =>
            -- reg_a = o3_X; reg_b = 2prime3; reg_acc = reg_o >> 256; o3_X = reg_o; operation : -s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_47 =>
            -- reg_a = o4_X; reg_b = 2prime4; reg_acc = reg_o >> 256; o4_X = reg_o; Enable sign a,b; operation : -s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_48 =>
            -- reg_a = o0_X; reg_b = 2prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '1';
            next_mac_sel_reg_s_reg_o_sign <= '1';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_49 =>
            -- reg_a = o1_X; reg_b = 2prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_50 =>
            -- reg_a = o2_X; reg_b = 2prime2; reg_acc = reg_o >> 256; o2_X = reg_o; operation : s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_51 =>
            -- reg_a = o3_X; reg_b = 2prime3; reg_acc = reg_o >> 256; o3_X = reg_o; operation : s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_52 =>
            -- reg_a = o4_X; reg_b = 2prime4; reg_acc = reg_o >> 256; o4_X = reg_o; Enable sign a,b; operation : s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_53 =>
            -- reg_a = o0_X; reg_b = 2prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '1';
            next_mac_sel_reg_s_reg_o_sign <= '1';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_54 =>
            -- reg_a = o1_X; reg_b = 2prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_55 =>
            -- reg_a = o2_X; reg_b = 2prime2; reg_acc = reg_o >> 256; o2_X = reg_o; operation : s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_56 =>
            -- reg_a = o3_X; reg_b = 2prime3; reg_acc = reg_o >> 256; o3_X = reg_o; operation : s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_57 =>
            -- reg_a = o4_X; reg_b = 2prime4; reg_acc = reg_o >> 256; o4_X = reg_o; Enable sign a,b; operation : s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_59 =>
            -- -- In case of size 6, 7, 8
            -- reg_a = a4_X; reg_b = b4_X; reg_acc = reg_o >> 256; o4_X = reg_o; operation : b +/- a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '1';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_60 =>
            -- -- In case of size 6
            -- reg_a = a5_X; reg_b = b5_X; reg_acc = reg_o >> 256; o5_X = reg_o; Enable sign a, b; operation : b +/- a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '1';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_61 =>
            -- reg_a = o0_X; reg_b = 2prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_positive; operation : -s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '1';
            next_mac_sel_reg_s_reg_o_sign <= '1';
            next_mac_reg_s_reg_o_positive <= '1';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_62 =>
            -- reg_a = o1_X; reg_b = 2prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : -s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_63 =>
            -- reg_a = o2_X; reg_b = 2prime2; reg_acc = reg_o >> 256; o2_X = reg_o; operation : -s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_64 =>
            -- reg_a = o3_X; reg_b = 2prime3; reg_acc = reg_o >> 256; o3_X = reg_o; operation : -s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_65 =>
            -- reg_a = o4_X; reg_b = 2prime4; reg_acc = reg_o >> 256; o4_X = reg_o; operation : -s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_66 =>
            -- reg_a = o5_X; reg_b = 2prime5; reg_acc = reg_o >> 256; o5_X = reg_o; Enable sign a,b; operation : -s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_67 =>
            -- reg_a = o0_X; reg_b = 2prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '1';
            next_mac_sel_reg_s_reg_o_sign <= '1';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_68 =>
            -- reg_a = o1_X; reg_b = 2prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_69 =>
            -- reg_a = o2_X; reg_b = 2prime2; reg_acc = reg_o >> 256; o2_X = reg_o; operation : s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_70 =>
            -- reg_a = o3_X; reg_b = 2prime3; reg_acc = reg_o >> 256; o3_X = reg_o; operation : s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_71 =>
            -- reg_a = o4_X; reg_b = 2prime4; reg_acc = reg_o >> 256; o4_X = reg_o; operation : s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_72 =>
            -- reg_a = o5_X; reg_b = 2prime5; reg_acc = reg_o >> 256; o5_X = reg_o; Enable sign a,b; operation : s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_73 =>
            -- reg_a = o0_X; reg_b = 2prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '1';
            next_mac_sel_reg_s_reg_o_sign <= '1';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_74 =>
            -- reg_a = o1_X; reg_b = 2prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_75 =>
            -- reg_a = o2_X; reg_b = 2prime2; reg_acc = reg_o >> 256; o2_X = reg_o; operation : s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_76 =>
            -- reg_a = o3_X; reg_b = 2prime3; reg_acc = reg_o >> 256; o3_X = reg_o; operation : s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_77 =>
            -- reg_a = o4_X; reg_b = 2prime4; reg_acc = reg_o >> 256; o4_X = reg_o; operation : s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_78 =>
            -- reg_a = o5_X; reg_b = 2prime5; reg_acc = reg_o >> 256; o5_X = reg_o; Enable sign a,b; operation : s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_80 =>
            -- -- In case of size 7, 8
            -- reg_a = a5_X; reg_b = b5_X; reg_acc = reg_o >> 256; o5_X = reg_o; operation : b +/- a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '1';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_81 =>
            -- -- In case of size 7
            -- reg_a = a6_X; reg_b = b6_X; reg_acc = reg_o >> 256; o6_X = reg_o; Enable sign a, b; operation : b +/- a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '1';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_82 =>
            -- reg_a = o0_X; reg_b = 2prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_positive; operation : -s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '1';
            next_mac_sel_reg_s_reg_o_sign <= '1';
            next_mac_reg_s_reg_o_positive <= '1';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_83 =>
            -- reg_a = o1_X; reg_b = 2prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : -s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_84 =>
            -- reg_a = o2_X; reg_b = 2prime2; reg_acc = reg_o >> 256; o2_X = reg_o; operation : -s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_85 =>
            -- reg_a = o3_X; reg_b = 2prime3; reg_acc = reg_o >> 256; o3_X = reg_o; operation : -s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_86 =>
            -- reg_a = o4_X; reg_b = 2prime4; reg_acc = reg_o >> 256; o4_X = reg_o; operation : -s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_87 =>
            -- reg_a = o5_X; reg_b = 2prime5; reg_acc = reg_o >> 256; o5_X = reg_o; operation : -s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_88 =>
            -- reg_a = o6_X; reg_b = 2prime6; reg_acc = reg_o >> 256; o6_X = reg_o; Enable sign a,b; operation : -s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_89 =>
            -- reg_a = o0_X; reg_b = 2prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '1';
            next_mac_sel_reg_s_reg_o_sign <= '1';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_90 =>
            -- reg_a = o1_X; reg_b = 2prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_91 =>
            -- reg_a = o2_X; reg_b = 2prime2; reg_acc = reg_o >> 256; o2_X = reg_o; operation : s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_92 =>
            -- reg_a = o3_X; reg_b = 2prime3; reg_acc = reg_o >> 256; o3_X = reg_o; operation : s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_93 =>
            -- reg_a = o4_X; reg_b = 2prime4; reg_acc = reg_o >> 256; o4_X = reg_o; operation : s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_94 =>
            -- reg_a = o5_X; reg_b = 2prime5; reg_acc = reg_o >> 256; o5_X = reg_o; operation : s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_95 =>
            -- reg_a = o6_X; reg_b = 2prime6; reg_acc = reg_o >> 256; o6_X = reg_o; Enable sign a,b; operation : s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_96 =>
            -- reg_a = o0_X; reg_b = 2prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '1';
            next_mac_sel_reg_s_reg_o_sign <= '1';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_97 =>
            -- reg_a = o1_X; reg_b = 2prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_98 =>
            -- reg_a = o2_X; reg_b = 2prime2; reg_acc = reg_o >> 256; o2_X = reg_o; operation : s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_99 =>
            -- reg_a = o3_X; reg_b = 2prime3; reg_acc = reg_o >> 256; o3_X = reg_o; operation : s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_100 =>
            -- reg_a = o4_X; reg_b = 2prime4; reg_acc = reg_o >> 256; o4_X = reg_o; operation : s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_101 =>
            -- reg_a = o5_X; reg_b = 2prime5; reg_acc = reg_o >> 256; o5_X = reg_o; operation : s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_102 =>
            -- reg_a = o6_X; reg_b = 2prime6; reg_acc = reg_o >> 256; o6_X = reg_o; Enable sign a,b; operation : s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_104 =>
            -- -- In case of size 8
            -- reg_a = a6_X; reg_b = b6_X; reg_acc = reg_o >> 256; o6_X = reg_o; operation : b +/- a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '1';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_105 =>
            -- reg_a = a7_X; reg_b = b7_X; reg_acc = reg_o >> 256; o7_X = reg_o; Enable sign a,b; operation : b +/- a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "111";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '1';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_106 =>
            -- reg_a = o0_X; reg_b = 2prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_positive; operation : -s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '1';
            next_mac_sel_reg_s_reg_o_sign <= '1';
            next_mac_reg_s_reg_o_positive <= '1';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_107 =>
            -- reg_a = o1_X; reg_b = 2prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : -s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_108 =>
            -- reg_a = o2_X; reg_b = 2prime2; reg_acc = reg_o >> 256; o2_X = reg_o; operation : -s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_109 =>
            -- reg_a = o3_X; reg_b = 2prime3; reg_acc = reg_o >> 256; o3_X = reg_o; operation : -s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_110 =>
            -- reg_a = o4_X; reg_b = 2prime4; reg_acc = reg_o >> 256; o4_X = reg_o; operation : -s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_111 =>
            -- reg_a = o5_X; reg_b = 2prime5; reg_acc = reg_o >> 256; o5_X = reg_o; operation : -s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_112 =>
            -- reg_a = o6_X; reg_b = 2prime6; reg_acc = reg_o >> 256; o6_X = reg_o; operation : -s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_113 =>
            -- reg_a = o7_X; reg_b = 2prime7; reg_acc = reg_o >> 256; o7_X = reg_o; Enable sign a,b; operation : -s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "111";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_114 =>
            -- reg_a = o0_X; reg_b = 2prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '1';
            next_mac_sel_reg_s_reg_o_sign <= '1';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_115 =>
            -- reg_a = o1_X; reg_b = 2prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_116 =>
            -- reg_a = o2_X; reg_b = 2prime2; reg_acc = reg_o >> 256; o2_X = reg_o; operation : s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_117 =>
            -- reg_a = o3_X; reg_b = 2prime3; reg_acc = reg_o >> 256; o3_X = reg_o; operation : s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_118 =>
            -- reg_a = o4_X; reg_b = 2prime4; reg_acc = reg_o >> 256; o4_X = reg_o; operation : s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "01";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_119 =>
            -- reg_a = o5_X; reg_b = 2prime5; reg_acc = reg_o >> 256; o5_X = reg_o; operation : s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_120 =>
            -- reg_a = o6_X; reg_b = 2prime6; reg_acc = reg_o >> 256; o6_X = reg_o; operation : s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_121 =>
            -- reg_a = o7_X; reg_b = 2prime7; reg_acc = reg_o >> 256; o7_X = reg_o; Enable sign a,b; operation : s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "111";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_122 =>
            -- reg_a = o0_X; reg_b = 2prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '1';
            next_mac_sel_reg_s_reg_o_sign <= '1';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_123 =>
            -- reg_a = o1_X; reg_b = 2prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_124 =>
            -- reg_a = o2_X; reg_b = 2prime2; reg_acc = reg_o >> 256; o2_X = reg_o; operation : s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_125 =>
            -- reg_a = o3_X; reg_b = 2prime3; reg_acc = reg_o >> 256; o3_X = reg_o; operation : s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_126 =>
            -- reg_a = o4_X; reg_b = 2prime4; reg_acc = reg_o >> 256; o4_X = reg_o; operation : s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_127 =>
            -- reg_a = o5_X; reg_b = 2prime5; reg_acc = reg_o >> 256; o5_X = reg_o; operation : s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_128 =>
            -- reg_a = o6_X; reg_b = 2prime6; reg_acc = reg_o >> 256; o6_X = reg_o; operation : s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_129 =>
            -- reg_a = o7_X; reg_b = 2prime7; reg_acc = reg_o >> 256; o7_X = reg_o; Enable sign a,b; operation : s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "01";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "111";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when nop_4_stages =>
        -- reg_a = 0; reg_b = 0; reg_acc = 0; operation : b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "11";
            next_mac_clear_reg_b <= '1';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when nop_8_stages =>
        -- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "11";
            next_mac_clear_reg_b <= '1';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
--        when others => 
--            next_sm_free_flag <= '0';
--            next_sm_rotation_size <= "11";
--            next_sm_circular_shift_enable <= '0';
--            next_sel_address_a <= '0';
--            next_sel_address_b_prime <= "00";
--            next_sm_specific_mac_address_a <= "000";
--            next_sm_specific_mac_address_b <= "000";
--            next_sm_specific_mac_address_o <= "000";
--            next_sm_specific_mac_next_address_o <= "001";
--            next_mac_enable_signed_a <= '0';
--            next_mac_enable_signed_b <= '0';
--            next_mac_sel_load_reg_a <= "11";
--            next_mac_clear_reg_b <= '1';
--            next_mac_clear_reg_acc <= '1';
--            next_mac_sel_shift_reg_o <= '0';
--            next_mac_enable_update_reg_s <= '0';
--            next_mac_sel_reg_s_reg_o_sign <= '0';
--            next_mac_reg_s_reg_o_positive <= '0';
--            next_sm_sign_a_mode <= '0';
--            next_sm_mac_operation_mode <= "10";
--            next_mac_enable_reg_s_mask <= '0';
--            next_mac_subtraction_reg_a_b <= '0';
--            next_mac_sel_multiply_two_a_b <= '0';
--            next_mac_sel_reg_y_output <= '0';
--            next_sm_mac_write_enable_output <= '0';
--            next_mac_memory_double_mode <= '0';
--            next_mac_memory_only_write_mode <= '0';
--            next_base_address_generator_o_increment_previous_address <= '0';
    end case;
end process;

update_state : process(actual_state, instruction_values_valid, instruction_type, prime_line_equal_one, operands_size, ultimate_operation)
begin
case (actual_state) is
        when reset =>
            next_state <= decode_instruction;
        when decode_instruction =>
            next_state <= decode_instruction;
            if(instruction_values_valid = '1') then
                if(instruction_type = "0000") then
                    if(operands_size = "000") then
                        next_state <= multiplication_direct_0;
                    else
                        next_state <= multiplication_direct_2;
                    end if;
                elsif(instruction_type = "0001") then
                    if(operands_size = "000") then
                        next_state <= square_direct_0;
                    else
                        next_state <= square_direct_2;
                    end if;
                elsif(instruction_type = "0010") then
                    case (prime_line_equal_one) is
                        when "00" =>
                            if(operands_size = "000") then
                                next_state <= multiplication_with_reduction_0;
                            else
                                next_state <= multiplication_with_reduction_5;
                            end if;
                        when "01" =>
                            if(operands_size = "000") then
                                next_state <= multiplication_with_reduction_special_prime_1_0;
                            else
                                next_state <= multiplication_with_reduction_special_prime_1_3;
                            end if;
                        when "10" =>
                            next_state <= multiplication_with_reduction_special_prime_2_0;
                        when "11" =>
                            next_state <= multiplication_with_reduction_special_prime_3_0;
                        when others =>
                            next_state <= decode_instruction;
                    end case;
                elsif(instruction_type = "0011") then
                    case (prime_line_equal_one) is
                        when "00" =>
                            if(operands_size = "000") then
                                next_state <= square_with_reduction_0;
                            else
                                next_state <= square_with_reduction_5;
                            end if;
                        when "01" =>
                            if(operands_size = "000") then
                                next_state <= square_with_reduction_special_prime_1_0;
                            else
                                next_state <= square_with_reduction_special_prime_1_3;
                            end if;
                        when "10" =>
                            next_state <= square_with_reduction_special_prime_2_0;
                        when "11" =>
                            next_state <= square_with_reduction_special_prime_3_0;
                        when others =>
                            next_state <= decode_instruction;
                    end case;
                elsif(instruction_type = "0100") then
                    if(operands_size = "000") then
                        next_state <= addition_subtraction_direct_0;
                    else
                        next_state <= addition_subtraction_direct_2;
                    end if;
                elsif(instruction_type = "0101") then
                    if(operands_size = "000") then
                        next_state <= iterative_modular_reduction_0;
                    elsif(operands_size = "001") then
                        next_state <= iterative_modular_reduction_5;
                    elsif(operands_size = "010") then
                        next_state <= iterative_modular_reduction_13;
                    elsif(operands_size = "011") then
                        next_state <= iterative_modular_reduction_24;
                    elsif(operands_size = "100") then
                        next_state <= iterative_modular_reduction_38;
                    elsif(operands_size = "101") then
                        next_state <= iterative_modular_reduction_55;
                    elsif(operands_size = "110") then
                        next_state <= iterative_modular_reduction_75;
                    else
                        next_state <= iterative_modular_reduction_98;
                    end if;
                elsif(instruction_type = "0110") then
                    if(operands_size = "000") then
                        next_state <= addition_subtraction_with_reduction_0;
                    else
                        next_state <= addition_subtraction_with_reduction_5;
                    end if;
                end if;
            end if;
        when multiplication_direct_0 =>
            next_state <= multiplication_direct_0;
            if(ultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when multiplication_direct_2 =>
            next_state <= multiplication_direct_2;
            if(ultimate_operation = '1') then
                if(operands_size = "001") then
                    next_state <= multiplication_direct_3;
                else
                    next_state <= multiplication_direct_7;
                end if;
            end if;
        when multiplication_direct_3 =>
            next_state <= multiplication_direct_3;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_4;
            end if;
        when multiplication_direct_4 =>
            next_state <= multiplication_direct_4;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_5;
            end if;
        when multiplication_direct_5 =>
            next_state <= multiplication_direct_5;
            if(ultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when multiplication_direct_7 =>
            next_state <= multiplication_direct_7;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_8;
            end if;
        when multiplication_direct_8 =>
            next_state <= multiplication_direct_8;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_9;
            end if;
        when multiplication_direct_9 =>
            next_state <= multiplication_direct_9;
            if(ultimate_operation = '1') then
                if(operands_size = "010") then
                    next_state <= multiplication_direct_10;
                else
                    next_state <= multiplication_direct_16;
                end if;
            end if;
        when multiplication_direct_10 =>
            next_state <= multiplication_direct_10;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_11;
            end if;
        when multiplication_direct_11 =>
            next_state <= multiplication_direct_11;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_12;
            end if;
        when multiplication_direct_12 =>
            next_state <= multiplication_direct_12;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_13;
            end if;
        when multiplication_direct_13 =>
            next_state <= multiplication_direct_13;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_14;
            end if;
        when multiplication_direct_14 =>
            next_state <= multiplication_direct_14;
            if(ultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when multiplication_direct_16 =>
            next_state <= multiplication_direct_16;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_17;
            end if;
        when multiplication_direct_17 =>
            next_state <= multiplication_direct_17;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_18;
            end if;
        when multiplication_direct_18 =>
            next_state <= multiplication_direct_18;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_19;
            end if;
        when multiplication_direct_19 =>
            next_state <= multiplication_direct_19;
            if(ultimate_operation = '1') then
                if(operands_size = "011") then
                    next_state <= multiplication_direct_20;
                else
                    next_state <= multiplication_direct_29;
                end if;
            end if;
        when multiplication_direct_20 =>
            next_state <= multiplication_direct_20;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_21;
            end if;
        when multiplication_direct_21 =>
            next_state <= multiplication_direct_21;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_22;
            end if;
        when multiplication_direct_22 =>
            next_state <= multiplication_direct_22;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_23;
            end if;
        when multiplication_direct_23 =>
            next_state <= multiplication_direct_23;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_24;
            end if;
        when multiplication_direct_24 =>
            next_state <= multiplication_direct_24;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_25;
            end if;
        when multiplication_direct_25 =>
            next_state <= multiplication_direct_25;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_26;
            end if;
        when multiplication_direct_26 =>
            next_state <= multiplication_direct_26;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_27;
            end if;
        when multiplication_direct_27 =>
            next_state <= multiplication_direct_27;
            if(ultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when multiplication_direct_29 =>
            next_state <= multiplication_direct_29;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_30;
            end if;
        when multiplication_direct_30 =>
            next_state <= multiplication_direct_30;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_31;
            end if;
        when multiplication_direct_31 =>
            next_state <= multiplication_direct_31;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_32;
            end if;
        when multiplication_direct_32 =>
            next_state <= multiplication_direct_32;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_33;
            end if;
        when multiplication_direct_33 =>
            next_state <= multiplication_direct_33;
            if(ultimate_operation = '1') then
                if(operands_size = "100") then
                    next_state <= multiplication_direct_34;
                else
                    next_state <= multiplication_direct_47;
                end if;
            end if;
        when multiplication_direct_34 =>
            next_state <= multiplication_direct_34;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_35;
            end if;
        when multiplication_direct_35 =>
            next_state <= multiplication_direct_35;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_36;
            end if;
        when multiplication_direct_36 =>
            next_state <= multiplication_direct_36;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_37;
            end if;
        when multiplication_direct_37 =>
            next_state <= multiplication_direct_37;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_38;
            end if;
        when multiplication_direct_38 =>
            next_state <= multiplication_direct_38;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_39;
            end if;
        when multiplication_direct_39 =>
            next_state <= multiplication_direct_39;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_40;
            end if;
        when multiplication_direct_40 =>
            next_state <= multiplication_direct_40;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_41;
            end if;
        when multiplication_direct_41 =>
            next_state <= multiplication_direct_41;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_42;
            end if;
        when multiplication_direct_42 =>
            next_state <= multiplication_direct_42;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_43;
            end if;
        when multiplication_direct_43 =>
            next_state <= multiplication_direct_43;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_44;
            end if;
        when multiplication_direct_44 =>
            next_state <= multiplication_direct_44;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_45;
            end if;
        when multiplication_direct_45 =>
            next_state <= multiplication_direct_45;
            if(ultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when multiplication_direct_47 =>
            next_state <= multiplication_direct_47;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_48;
            end if;
        when multiplication_direct_48 =>
            next_state <= multiplication_direct_48;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_49;
            end if;
        when multiplication_direct_49 =>
            next_state <= multiplication_direct_49;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_50;
            end if;
        when multiplication_direct_50 =>
            next_state <= multiplication_direct_50;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_51;
            end if;
        when multiplication_direct_51 =>
            next_state <= multiplication_direct_51;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_52;
            end if;
        when multiplication_direct_52 =>
            next_state <= multiplication_direct_52;
            if(ultimate_operation = '1') then
                if(operands_size = "101") then
                    next_state <= multiplication_direct_53;
                else
                    next_state <= multiplication_direct_71;
                end if;
            end if;
        when multiplication_direct_53 =>
            next_state <= multiplication_direct_53;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_54;
            end if;
        when multiplication_direct_54 =>
            next_state <= multiplication_direct_54;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_55;
            end if;
        when multiplication_direct_55 =>
            next_state <= multiplication_direct_55;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_56;
            end if;
        when multiplication_direct_56 =>
            next_state <= multiplication_direct_56;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_57;
            end if;
        when multiplication_direct_57 =>
            next_state <= multiplication_direct_57;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_58;
            end if;
        when multiplication_direct_58 =>
            next_state <= multiplication_direct_58;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_59;
            end if;
        when multiplication_direct_59 =>
            next_state <= multiplication_direct_59;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_60;
            end if;
        when multiplication_direct_60 =>
            next_state <= multiplication_direct_60;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_61;
            end if;
        when multiplication_direct_61 =>
            next_state <= multiplication_direct_61;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_62;
            end if;
        when multiplication_direct_62 =>
            next_state <= multiplication_direct_62;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_63;
            end if;
        when multiplication_direct_63 =>
            next_state <= multiplication_direct_63;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_64;
            end if;
        when multiplication_direct_64 =>
            next_state <= multiplication_direct_64;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_65;
            end if;
        when multiplication_direct_65 =>
            next_state <= multiplication_direct_65;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_66;
            end if;
        when multiplication_direct_66 =>
            next_state <= multiplication_direct_66;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_67;
            end if;
        when multiplication_direct_67 =>
            next_state <= multiplication_direct_67;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_68;
            end if;
        when multiplication_direct_68 =>
            next_state <= multiplication_direct_68;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_69;
            end if;
        when multiplication_direct_69 =>
            next_state <= multiplication_direct_69;
            if(ultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when multiplication_direct_71 =>
            next_state <= multiplication_direct_71;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_72;
            end if;
        when multiplication_direct_72 =>
            next_state <= multiplication_direct_72;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_73;
            end if;
        when multiplication_direct_73 =>
            next_state <= multiplication_direct_73;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_74;
            end if;
        when multiplication_direct_74 =>
            next_state <= multiplication_direct_74;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_75;
            end if;
        when multiplication_direct_75 =>
            next_state <= multiplication_direct_75;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_76;
            end if;
        when multiplication_direct_76 =>
            next_state <= multiplication_direct_76;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_77;
            end if;
        when multiplication_direct_77 =>
            next_state <= multiplication_direct_77;
            if(ultimate_operation = '1') then
                if(operands_size = "110") then
                    next_state <= multiplication_direct_78;
                else
                    next_state <= multiplication_direct_102;
                end if;
            end if;
        when multiplication_direct_78 =>
            next_state <= multiplication_direct_78;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_79;
            end if;
        when multiplication_direct_79 =>
            next_state <= multiplication_direct_79;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_80;
            end if;
        when multiplication_direct_80 =>
            next_state <= multiplication_direct_80;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_81;
            end if;
        when multiplication_direct_81 =>
            next_state <= multiplication_direct_81;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_82;
            end if;
        when multiplication_direct_82 =>
            next_state <= multiplication_direct_82;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_83;
            end if;
        when multiplication_direct_83 =>
            next_state <= multiplication_direct_83;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_84;
            end if;
        when multiplication_direct_84 =>
            next_state <= multiplication_direct_84;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_85;
            end if;
        when multiplication_direct_85 =>
            next_state <= multiplication_direct_85;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_86;
            end if;
        when multiplication_direct_86 =>
            next_state <= multiplication_direct_86;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_87;
            end if;
        when multiplication_direct_87 =>
            next_state <= multiplication_direct_87;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_88;
            end if;
        when multiplication_direct_88 =>
            next_state <= multiplication_direct_88;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_89;
            end if;
        when multiplication_direct_89 =>
            next_state <= multiplication_direct_89;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_90;
            end if;
        when multiplication_direct_90 =>
            next_state <= multiplication_direct_90;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_91;
            end if;
        when multiplication_direct_91 =>
            next_state <= multiplication_direct_91;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_92;
            end if;
        when multiplication_direct_92 =>
            next_state <= multiplication_direct_92;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_93;
            end if;
        when multiplication_direct_93 =>
            next_state <= multiplication_direct_93;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_94;
            end if;
        when multiplication_direct_94 =>
            next_state <= multiplication_direct_94;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_95;
            end if;
        when multiplication_direct_95 =>
            next_state <= multiplication_direct_95;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_96;
            end if;
        when multiplication_direct_96 =>
            next_state <= multiplication_direct_96;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_97;
            end if;
        when multiplication_direct_97 =>
            next_state <= multiplication_direct_97;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_98;
            end if;
        when multiplication_direct_98 =>
            next_state <= multiplication_direct_98;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_99;
            end if;
        when multiplication_direct_99 =>
            next_state <= multiplication_direct_99;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_100;
            end if;
        when multiplication_direct_100 =>
            next_state <= multiplication_direct_100;
            if(ultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when multiplication_direct_102 =>
            next_state <= multiplication_direct_102;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_103;
            end if;
        when multiplication_direct_103 =>
            next_state <= multiplication_direct_103;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_104;
            end if;
        when multiplication_direct_104 =>
            next_state <= multiplication_direct_104;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_105;
            end if;
        when multiplication_direct_105 =>
            next_state <= multiplication_direct_105;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_106;
            end if;
        when multiplication_direct_106 =>
            next_state <= multiplication_direct_106;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_107;
            end if;
        when multiplication_direct_107 =>
            next_state <= multiplication_direct_107;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_108;
            end if;
        when multiplication_direct_108 =>
            next_state <= multiplication_direct_108;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_109;
            end if;
        when multiplication_direct_109 =>
            next_state <= multiplication_direct_109;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_110;
            end if;
        when multiplication_direct_110 =>
            next_state <= multiplication_direct_110;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_111;
            end if;
        when multiplication_direct_111 =>
            next_state <= multiplication_direct_111;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_112;
            end if;
        when multiplication_direct_112 =>
            next_state <= multiplication_direct_112;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_113;
            end if;
        when multiplication_direct_113 =>
            next_state <= multiplication_direct_113;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_114;
            end if;
        when multiplication_direct_114 =>
            next_state <= multiplication_direct_114;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_115;
            end if;
        when multiplication_direct_115 =>
            next_state <= multiplication_direct_115;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_116;
            end if;
        when multiplication_direct_116 =>
            next_state <= multiplication_direct_116;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_117;
            end if;
        when multiplication_direct_117 =>
            next_state <= multiplication_direct_117;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_118;
            end if;
        when multiplication_direct_118 =>
            next_state <= multiplication_direct_118;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_119;
            end if;
        when multiplication_direct_119 =>
            next_state <= multiplication_direct_119;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_120;
            end if;
        when multiplication_direct_120 =>
            next_state <= multiplication_direct_120;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_121;
            end if;
        when multiplication_direct_121 =>
            next_state <= multiplication_direct_121;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_122;
            end if;
        when multiplication_direct_122 =>
            next_state <= multiplication_direct_122;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_123;
            end if;
        when multiplication_direct_123 =>
            next_state <= multiplication_direct_123;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_124;
            end if;
        when multiplication_direct_124 =>
            next_state <= multiplication_direct_124;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_125;
            end if;
        when multiplication_direct_125 =>
            next_state <= multiplication_direct_125;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_126;
            end if;
        when multiplication_direct_126 =>
            next_state <= multiplication_direct_126;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_127;
            end if;
        when multiplication_direct_127 =>
            next_state <= multiplication_direct_127;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_128;
            end if;
        when multiplication_direct_128 =>
            next_state <= multiplication_direct_128;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_129;
            end if;
        when multiplication_direct_129 =>
            next_state <= multiplication_direct_129;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_130;
            end if;
        when multiplication_direct_130 =>
            next_state <= multiplication_direct_130;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_131;
            end if;
        when multiplication_direct_131 =>
            next_state <= multiplication_direct_131;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_132;
            end if;
        when multiplication_direct_132 =>
            next_state <= multiplication_direct_132;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_133;
            end if;
        when multiplication_direct_133 =>
            next_state <= multiplication_direct_133;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_134;
            end if;
        when multiplication_direct_134 =>
            next_state <= multiplication_direct_134;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_135;
            end if;
        when multiplication_direct_135 =>
            next_state <= multiplication_direct_135;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_136;
            end if;
        when multiplication_direct_136 =>
            next_state <= multiplication_direct_136;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_137;
            end if;
        when multiplication_direct_137 =>
            next_state <= multiplication_direct_137;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_138;
            end if;
        when multiplication_direct_138 =>
            next_state <= multiplication_direct_138;
            if(ultimate_operation = '1') then
                next_state <= multiplication_direct_139;
            end if;
        when multiplication_direct_139 =>
            next_state <= multiplication_direct_139;
            if(ultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when square_direct_0 => 
            next_state <= square_direct_0;
            if(ultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when square_direct_2 => 
            next_state <= square_direct_2;
            if(ultimate_operation = '1') then
                if(operands_size = "001") then
                    next_state <= square_direct_3;
                else
                    next_state <= square_direct_6;
                end if;
            end if;
        when square_direct_3 => 
            next_state <= square_direct_3;
            if(ultimate_operation = '1') then
                next_state <= square_direct_4;
            end if;
        when square_direct_4 => 
            next_state <= square_direct_4;
            if(ultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when square_direct_6 => 
            next_state <= square_direct_6;
            if(ultimate_operation = '1') then
                next_state <= square_direct_7;
            end if;
        when square_direct_7 => 
            next_state <= square_direct_7;
            if(ultimate_operation = '1') then
                if(operands_size = "010") then
                    next_state <= square_direct_8;
                else
                    next_state <= square_direct_12;
                end if;
            end if;
        when square_direct_8 => 
            next_state <= square_direct_8;
            if(ultimate_operation = '1') then
                next_state <= square_direct_9;
            end if;
        when square_direct_9 => 
            next_state <= square_direct_9;
            if(ultimate_operation = '1') then
                next_state <= square_direct_10;
            end if;
        when square_direct_10 => 
            next_state <= square_direct_10;
            if(ultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when square_direct_12 => 
            next_state <= square_direct_12;
            if(ultimate_operation = '1') then
                next_state <= square_direct_13;
            end if;
        when square_direct_13 => 
            next_state <= square_direct_13;
            if(ultimate_operation = '1') then
                if(operands_size = "011") then
                    next_state <= square_direct_14;
                else
                    next_state <= square_direct_20;
                end if;
            end if;
        when square_direct_14 => 
            next_state <= square_direct_14;
            if(ultimate_operation = '1') then
                next_state <= square_direct_15;
            end if;
        when square_direct_15 => 
            next_state <= square_direct_15;
            if(ultimate_operation = '1') then
                next_state <= square_direct_16;
            end if;
        when square_direct_16 => 
            next_state <= square_direct_16;
            if(ultimate_operation = '1') then
                next_state <= square_direct_17;
            end if;
        when square_direct_17 => 
            next_state <= square_direct_17;
            if(ultimate_operation = '1') then
                next_state <= square_direct_18;
            end if;
        when square_direct_18 => 
            next_state <= square_direct_18;
            if(ultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when square_direct_20 => 
            next_state <= square_direct_20;
            if(ultimate_operation = '1') then
                next_state <= square_direct_21;
            end if;
        when square_direct_21 => 
            next_state <= square_direct_21;
            if(ultimate_operation = '1') then
                next_state <= square_direct_22;
            end if;
        when square_direct_22 => 
            next_state <= square_direct_22;
            if(ultimate_operation = '1') then
                if(operands_size = "100") then
                    next_state <= square_direct_23;
                else
                    next_state <= square_direct_31;
                end if;
            end if;
        when square_direct_23 => 
            next_state <= square_direct_23;
            if(ultimate_operation = '1') then
                next_state <= square_direct_24;
            end if;
        when square_direct_24 => 
            next_state <= square_direct_24;
            if(ultimate_operation = '1') then
                next_state <= square_direct_25;
            end if;
        when square_direct_25 => 
            next_state <= square_direct_25;
            if(ultimate_operation = '1') then
                next_state <= square_direct_26;
            end if;
        when square_direct_26 => 
            next_state <= square_direct_26;
            if(ultimate_operation = '1') then
                next_state <= square_direct_27;
            end if;
        when square_direct_27 => 
            next_state <= square_direct_27;
            if(ultimate_operation = '1') then
                next_state <= square_direct_28;
            end if;
        when square_direct_28 => 
            next_state <= square_direct_28;
            if(ultimate_operation = '1') then
                next_state <= square_direct_29;
            end if;
        when square_direct_29 => 
            next_state <= square_direct_29;
            if(ultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when square_direct_31 => 
            next_state <= square_direct_31;
            if(ultimate_operation = '1') then
                next_state <= square_direct_32;
            end if;
        when square_direct_32 => 
            next_state <= square_direct_32;
            if(ultimate_operation = '1') then
                next_state <= square_direct_33;
            end if;
        when square_direct_33 => 
            next_state <= square_direct_33;
            if(ultimate_operation = '1') then
                if(operands_size = "101") then
                    next_state <= square_direct_34;
                else
                    next_state <= square_direct_45;
                end if;
            end if;
        when square_direct_34 => 
            next_state <= square_direct_34;
            if(ultimate_operation = '1') then
                next_state <= square_direct_35;
            end if;
        when square_direct_35 => 
            next_state <= square_direct_35;
            if(ultimate_operation = '1') then
                next_state <= square_direct_36;
            end if;
        when square_direct_36 => 
            next_state <= square_direct_36;
            if(ultimate_operation = '1') then
                next_state <= square_direct_37;
            end if;
        when square_direct_37 => 
            next_state <= square_direct_37;
            if(ultimate_operation = '1') then
                next_state <= square_direct_38;
            end if;
        when square_direct_38 => 
            next_state <= square_direct_38;
            if(ultimate_operation = '1') then
                next_state <= square_direct_39;
            end if;
        when square_direct_39 => 
            next_state <= square_direct_39;
            if(ultimate_operation = '1') then
                next_state <= square_direct_40;
            end if;
        when square_direct_40 => 
            next_state <= square_direct_40;
            if(ultimate_operation = '1') then
                next_state <= square_direct_41;
            end if;
        when square_direct_41 => 
            next_state <= square_direct_41;
            if(ultimate_operation = '1') then
                next_state <= square_direct_42;
            end if;
        when square_direct_42 => 
            next_state <= square_direct_42;
            if(ultimate_operation = '1') then
                next_state <= square_direct_43;
            end if;
        when square_direct_43 => 
            next_state <= square_direct_43;
            if(ultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when square_direct_45 => 
            next_state <= square_direct_45;
            if(ultimate_operation = '1') then
                next_state <= square_direct_46;
            end if;
        when square_direct_46 => 
            next_state <= square_direct_46;
            if(ultimate_operation = '1') then
                next_state <= square_direct_47;
            end if;
        when square_direct_47 => 
            next_state <= square_direct_47;
            if(ultimate_operation = '1') then
                next_state <= square_direct_48;
            end if;
        when square_direct_48 => 
            next_state <= square_direct_48;
            if(ultimate_operation = '1') then
                if(operands_size = "110") then
                    next_state <= square_direct_49;
                else
                    next_state <= square_direct_63;
                end if;
            end if;
        when square_direct_49 => 
            next_state <= square_direct_49;
            if(ultimate_operation = '1') then
                next_state <= square_direct_50;
            end if;
        when square_direct_50 => 
            next_state <= square_direct_50;
            if(ultimate_operation = '1') then
                next_state <= square_direct_51;
            end if;
        when square_direct_51 => 
            next_state <= square_direct_51;
            if(ultimate_operation = '1') then
                next_state <= square_direct_52;
            end if;
        when square_direct_52 => 
            next_state <= square_direct_52;
            if(ultimate_operation = '1') then
                next_state <= square_direct_53;
            end if;
        when square_direct_53 => 
            next_state <= square_direct_53;
            if(ultimate_operation = '1') then
                next_state <= square_direct_54;
            end if;
        when square_direct_54 => 
            next_state <= square_direct_54;
            if(ultimate_operation = '1') then
                next_state <= square_direct_55;
            end if;
        when square_direct_55 => 
            next_state <= square_direct_55;
            if(ultimate_operation = '1') then
                next_state <= square_direct_56;
            end if;
        when square_direct_56 => 
            next_state <= square_direct_56;
            if(ultimate_operation = '1') then
                next_state <= square_direct_57;
            end if;
        when square_direct_57 => 
            next_state <= square_direct_57;
            if(ultimate_operation = '1') then
                next_state <= square_direct_58;
            end if;
        when square_direct_58 => 
            next_state <= square_direct_58;
            if(ultimate_operation = '1') then
                next_state <= square_direct_59;
            end if;
        when square_direct_59 => 
            next_state <= square_direct_59;
            if(ultimate_operation = '1') then
                next_state <= square_direct_60;
            end if;
        when square_direct_60 => 
            next_state <= square_direct_60;
            if(ultimate_operation = '1') then
                next_state <= square_direct_61;
            end if;
        when square_direct_61 => 
            next_state <= square_direct_61;
            if(ultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when square_direct_63 => 
            next_state <= square_direct_63;
            if(ultimate_operation = '1') then
                next_state <= square_direct_64;
            end if;
        when square_direct_64 => 
            next_state <= square_direct_64;
            if(ultimate_operation = '1') then
                next_state <= square_direct_65;
            end if;
        when square_direct_65 => 
            next_state <= square_direct_65;
            if(ultimate_operation = '1') then
                next_state <= square_direct_66;
            end if;
        when square_direct_66 => 
            next_state <= square_direct_66;
            if(ultimate_operation = '1') then
                next_state <= square_direct_67;
            end if;
        when square_direct_67 => 
            next_state <= square_direct_67;
            if(ultimate_operation = '1') then
                next_state <= square_direct_68;
            end if;
        when square_direct_68 => 
            next_state <= square_direct_68;
            if(ultimate_operation = '1') then
                next_state <= square_direct_69;
            end if;
        when square_direct_69 => 
            next_state <= square_direct_69;
            if(ultimate_operation = '1') then
                next_state <= square_direct_70;
            end if;
        when square_direct_70 => 
            next_state <= square_direct_70;
            if(ultimate_operation = '1') then
                next_state <= square_direct_71;
            end if;
        when square_direct_71 => 
            next_state <= square_direct_71;
            if(ultimate_operation = '1') then
                next_state <= square_direct_72;
            end if;
        when square_direct_72 => 
            next_state <= square_direct_72;
            if(ultimate_operation = '1') then
                next_state <= square_direct_73;
            end if;
        when square_direct_73 => 
            next_state <= square_direct_73;
            if(ultimate_operation = '1') then
                next_state <= square_direct_74;
            end if;
        when square_direct_74 => 
            next_state <= square_direct_74;
            if(ultimate_operation = '1') then
                next_state <= square_direct_75;
            end if;
        when square_direct_75 => 
            next_state <= square_direct_75;
            if(ultimate_operation = '1') then
                next_state <= square_direct_76;
            end if;
        when square_direct_76 => 
            next_state <= square_direct_76;
            if(ultimate_operation = '1') then
                next_state <= square_direct_77;
            end if;
        when square_direct_77 => 
            next_state <= square_direct_77;
            if(ultimate_operation = '1') then
                next_state <= square_direct_78;
            end if;
        when square_direct_78 => 
            next_state <= square_direct_78;
            if(ultimate_operation = '1') then
                next_state <= square_direct_79;
            end if;
        when square_direct_79 => 
            next_state <= square_direct_79;
            if(ultimate_operation = '1') then
                next_state <= square_direct_80;
            end if;
        when square_direct_80 => 
            next_state <= square_direct_80;
            if(ultimate_operation = '1') then
                next_state <= square_direct_81;
            end if;
        when square_direct_81 => 
            next_state <= square_direct_81;
            if(ultimate_operation = '1') then
                next_state <= square_direct_82;
            end if;
        when square_direct_82 => 
            next_state <= square_direct_82;
            if(ultimate_operation = '1') then
                next_state <= square_direct_83;
            end if;
        when square_direct_83 => 
            next_state <= square_direct_83;
            if(ultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when multiplication_with_reduction_0 => 
            next_state <= multiplication_with_reduction_0;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_1;
            end if;
        when multiplication_with_reduction_1 => 
            next_state <= multiplication_with_reduction_1;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_2;
            end if;
        when multiplication_with_reduction_2 => 
            next_state <= multiplication_with_reduction_2;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_3;
            end if;
        when multiplication_with_reduction_3 => 
            next_state <= multiplication_with_reduction_3;
            if(ultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when multiplication_with_reduction_5 => 
            next_state <= multiplication_with_reduction_5;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_6;
            end if;
        when multiplication_with_reduction_6 => 
            next_state <= multiplication_with_reduction_6;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_7;
            end if;
        when multiplication_with_reduction_7 => 
            next_state <= multiplication_with_reduction_7;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_8;
            end if;
        when multiplication_with_reduction_8 => 
            next_state <= multiplication_with_reduction_8;
            if(ultimate_operation = '1') then
                if(operands_size = "001") then
                    next_state <= multiplication_with_reduction_9;
                else
                    next_state <= multiplication_with_reduction_16;
                end if;
            end if;
        when multiplication_with_reduction_9 => 
            next_state <= multiplication_with_reduction_9;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_10;
            end if;
        when multiplication_with_reduction_10 => 
            next_state <= multiplication_with_reduction_10;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_11;
            end if;
        when multiplication_with_reduction_11 => 
            next_state <= multiplication_with_reduction_11;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_12;
            end if;
        when multiplication_with_reduction_12 => 
            next_state <= multiplication_with_reduction_12;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_13;
            end if;
        when multiplication_with_reduction_13 => 
            next_state <= multiplication_with_reduction_13;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_14;
            end if;
        when multiplication_with_reduction_14 => 
            next_state <= multiplication_with_reduction_14;
            if(ultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when multiplication_with_reduction_16 => 
            next_state <= multiplication_with_reduction_16;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_17;
            end if;
        when multiplication_with_reduction_17 => 
            next_state <= multiplication_with_reduction_17;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_18;
            end if;
        when multiplication_with_reduction_18 => 
            next_state <= multiplication_with_reduction_18;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_19;
            end if;
        when multiplication_with_reduction_19 => 
            next_state <= multiplication_with_reduction_19;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_20;
            end if;
        when multiplication_with_reduction_20 => 
            next_state <= multiplication_with_reduction_20;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_21;
            end if;
        when multiplication_with_reduction_21 => 
            next_state <= multiplication_with_reduction_21;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_22;
            end if;
        when multiplication_with_reduction_22 => 
            next_state <= multiplication_with_reduction_22;
            if(ultimate_operation = '1') then
                if(operands_size = "010") then
                    next_state <= multiplication_with_reduction_23;
                else
                    next_state <= multiplication_with_reduction_34;
                end if;
            end if;
        when multiplication_with_reduction_23 => 
            next_state <= multiplication_with_reduction_23;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_24;
            end if;
        when multiplication_with_reduction_24 => 
            next_state <= multiplication_with_reduction_24;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_25;
            end if;
        when multiplication_with_reduction_25 => 
            next_state <= multiplication_with_reduction_25;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_26;
            end if;
        when multiplication_with_reduction_26 => 
            next_state <= multiplication_with_reduction_26;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_27;
            end if;
        when multiplication_with_reduction_27 => 
            next_state <= multiplication_with_reduction_27;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_28;
            end if;
        when multiplication_with_reduction_28 => 
            next_state <= multiplication_with_reduction_28;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_29;
            end if;
        when multiplication_with_reduction_29 => 
            next_state <= multiplication_with_reduction_29;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_30;
            end if;
        when multiplication_with_reduction_30 => 
            next_state <= multiplication_with_reduction_30;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_31;
            end if;
        when multiplication_with_reduction_31 => 
            next_state <= multiplication_with_reduction_31;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_32;
            end if;
        when multiplication_with_reduction_32 => 
            next_state <= multiplication_with_reduction_32;
            if(ultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when multiplication_with_reduction_34 => 
            next_state <= multiplication_with_reduction_34;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_35;
            end if;
        when multiplication_with_reduction_35 => 
            next_state <= multiplication_with_reduction_35;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_36;
            end if;
        when multiplication_with_reduction_36 => 
            next_state <= multiplication_with_reduction_36;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_37;
            end if;
        when multiplication_with_reduction_37 => 
            next_state <= multiplication_with_reduction_37;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_38;
            end if;
        when multiplication_with_reduction_38 => 
            next_state <= multiplication_with_reduction_38;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_39;
            end if;
        when multiplication_with_reduction_39 => 
            next_state <= multiplication_with_reduction_39;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_40;
            end if;
        when multiplication_with_reduction_40 => 
            next_state <= multiplication_with_reduction_40;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_41;
            end if;
        when multiplication_with_reduction_41 => 
            next_state <= multiplication_with_reduction_41;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_42;
            end if;
        when multiplication_with_reduction_42 => 
            next_state <= multiplication_with_reduction_42;
            if(ultimate_operation = '1') then
                if(operands_size = "011") then
                    next_state <= multiplication_with_reduction_43;
                else
                    next_state <= multiplication_with_reduction_60;
                end if;
            end if;
        when multiplication_with_reduction_43 => 
            next_state <= multiplication_with_reduction_43;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_44;
            end if;
        when multiplication_with_reduction_44 => 
            next_state <= multiplication_with_reduction_44;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_45;
            end if;
        when multiplication_with_reduction_45 => 
            next_state <= multiplication_with_reduction_45;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_46;
            end if;
        when multiplication_with_reduction_46 => 
            next_state <= multiplication_with_reduction_46;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_47;
            end if;
        when multiplication_with_reduction_47 => 
            next_state <= multiplication_with_reduction_47;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_48;
            end if;
        when multiplication_with_reduction_48 => 
            next_state <= multiplication_with_reduction_48;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_49;
            end if;
        when multiplication_with_reduction_49 => 
            next_state <= multiplication_with_reduction_49;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_50;
            end if;
        when multiplication_with_reduction_50 => 
            next_state <= multiplication_with_reduction_50;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_51;
            end if;
        when multiplication_with_reduction_51 => 
            next_state <= multiplication_with_reduction_51;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_52;
            end if;
        when multiplication_with_reduction_52 => 
            next_state <= multiplication_with_reduction_52;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_53;
            end if;
        when multiplication_with_reduction_53 => 
            next_state <= multiplication_with_reduction_53;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_54;
            end if;
        when multiplication_with_reduction_54 => 
            next_state <= multiplication_with_reduction_54;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_55;
            end if;
        when multiplication_with_reduction_55 => 
            next_state <= multiplication_with_reduction_55;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_56;
            end if;
        when multiplication_with_reduction_56 => 
            next_state <= multiplication_with_reduction_56;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_57;
            end if;
        when multiplication_with_reduction_57 => 
            next_state <= multiplication_with_reduction_57;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_58;
            end if;
        when multiplication_with_reduction_58 => 
            next_state <= multiplication_with_reduction_58;
            if(ultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when multiplication_with_reduction_60 => 
            next_state <= multiplication_with_reduction_60;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_61;
            end if;
        when multiplication_with_reduction_61 => 
            next_state <= multiplication_with_reduction_61;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_62;
            end if;
        when multiplication_with_reduction_62 => 
            next_state <= multiplication_with_reduction_62;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_63;
            end if;
        when multiplication_with_reduction_63 => 
            next_state <= multiplication_with_reduction_63;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_64;
            end if;
        when multiplication_with_reduction_64 => 
            next_state <= multiplication_with_reduction_64;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_65;
            end if;
        when multiplication_with_reduction_65 => 
            next_state <= multiplication_with_reduction_65;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_66;
            end if;
        when multiplication_with_reduction_66 => 
            next_state <= multiplication_with_reduction_66;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_67;
            end if;
        when multiplication_with_reduction_67 => 
            next_state <= multiplication_with_reduction_67;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_68;
            end if;
        when multiplication_with_reduction_68 => 
            next_state <= multiplication_with_reduction_68;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_69;
            end if;
        when multiplication_with_reduction_69 => 
            next_state <= multiplication_with_reduction_69;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_70;
            end if;
        when multiplication_with_reduction_70 => 
            next_state <= multiplication_with_reduction_70;
            if(ultimate_operation = '1') then
                if(operands_size = "100") then
                    next_state <= multiplication_with_reduction_71;
                else
                    next_state <= multiplication_with_reduction_96;
                end if;
            end if;
        when multiplication_with_reduction_71 => 
            next_state <= multiplication_with_reduction_71;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_72;
            end if;
        when multiplication_with_reduction_72 => 
            next_state <= multiplication_with_reduction_72;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_73;
            end if;
        when multiplication_with_reduction_73 => 
            next_state <= multiplication_with_reduction_73;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_74;
            end if;
        when multiplication_with_reduction_74 => 
            next_state <= multiplication_with_reduction_74;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_75;
            end if;
        when multiplication_with_reduction_75 => 
            next_state <= multiplication_with_reduction_75;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_76;
            end if;
        when multiplication_with_reduction_76 => 
            next_state <= multiplication_with_reduction_76;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_77;
            end if;
        when multiplication_with_reduction_77 => 
            next_state <= multiplication_with_reduction_77;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_78;
            end if;
        when multiplication_with_reduction_78 => 
            next_state <= multiplication_with_reduction_78;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_79;
            end if;
        when multiplication_with_reduction_79 => 
            next_state <= multiplication_with_reduction_79;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_80;
            end if;
        when multiplication_with_reduction_80 => 
            next_state <= multiplication_with_reduction_80;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_81;
            end if;
        when multiplication_with_reduction_81 => 
            next_state <= multiplication_with_reduction_81;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_82;
            end if;
        when multiplication_with_reduction_82 => 
            next_state <= multiplication_with_reduction_82;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_83;
            end if;
        when multiplication_with_reduction_83 => 
            next_state <= multiplication_with_reduction_83;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_84;
            end if;
        when multiplication_with_reduction_84 => 
            next_state <= multiplication_with_reduction_84;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_85;
            end if;
        when multiplication_with_reduction_85 => 
            next_state <= multiplication_with_reduction_85;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_86;
            end if;
        when multiplication_with_reduction_86 => 
            next_state <= multiplication_with_reduction_86;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_87;
            end if;
        when multiplication_with_reduction_87 => 
            next_state <= multiplication_with_reduction_87;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_88;
            end if;
        when multiplication_with_reduction_88 => 
            next_state <= multiplication_with_reduction_88;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_89;
            end if;
        when multiplication_with_reduction_89 => 
            next_state <= multiplication_with_reduction_89;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_90;
            end if;
        when multiplication_with_reduction_90 => 
            next_state <= multiplication_with_reduction_90;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_91;
            end if;
        when multiplication_with_reduction_91 => 
            next_state <= multiplication_with_reduction_91;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_92;
            end if;
        when multiplication_with_reduction_92 => 
            next_state <= multiplication_with_reduction_92;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_93;
            end if;
        when multiplication_with_reduction_93 => 
            next_state <= multiplication_with_reduction_93;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_94;
            end if;
        when multiplication_with_reduction_94 => 
            next_state <= multiplication_with_reduction_94;
            if(ultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when multiplication_with_reduction_96 => 
            next_state <= multiplication_with_reduction_96;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_97;
            end if;
        when multiplication_with_reduction_97 => 
            next_state <= multiplication_with_reduction_97;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_98;
            end if;
        when multiplication_with_reduction_98 => 
            next_state <= multiplication_with_reduction_98;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_99;
            end if;
        when multiplication_with_reduction_99 => 
            next_state <= multiplication_with_reduction_99;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_100;
            end if;
        when multiplication_with_reduction_100 => 
            next_state <= multiplication_with_reduction_100;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_101;
            end if;
        when multiplication_with_reduction_101 => 
            next_state <= multiplication_with_reduction_101;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_102;
            end if;
        when multiplication_with_reduction_102 => 
            next_state <= multiplication_with_reduction_102;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_103;
            end if;
        when multiplication_with_reduction_103 => 
            next_state <= multiplication_with_reduction_103;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_104;
            end if;
        when multiplication_with_reduction_104 => 
            next_state <= multiplication_with_reduction_104;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_105;
            end if;
        when multiplication_with_reduction_105 => 
            next_state <= multiplication_with_reduction_105;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_106;
            end if;
        when multiplication_with_reduction_106 => 
            next_state <= multiplication_with_reduction_106;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_107;
            end if;
        when multiplication_with_reduction_107 => 
            next_state <= multiplication_with_reduction_107;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_108;
            end if;
        when multiplication_with_reduction_108 => 
            next_state <= multiplication_with_reduction_108;
            if(ultimate_operation = '1') then
                if(operands_size = "101") then
                    next_state <= multiplication_with_reduction_109;
                else
                    next_state <= multiplication_with_reduction_144;
                end if;
            end if;
        when multiplication_with_reduction_109 => 
            next_state <= multiplication_with_reduction_109;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_110;
            end if;
        when multiplication_with_reduction_110 => 
            next_state <= multiplication_with_reduction_110;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_111;
            end if;
        when multiplication_with_reduction_111 => 
            next_state <= multiplication_with_reduction_111;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_112;
            end if;
        when multiplication_with_reduction_112 => 
            next_state <= multiplication_with_reduction_112;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_113;
            end if;
        when multiplication_with_reduction_113 => 
            next_state <= multiplication_with_reduction_113;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_114;
            end if;
        when multiplication_with_reduction_114 => 
            next_state <= multiplication_with_reduction_114;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_115;
            end if;
        when multiplication_with_reduction_115 => 
            next_state <= multiplication_with_reduction_115;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_116;
            end if;
        when multiplication_with_reduction_116 => 
            next_state <= multiplication_with_reduction_116;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_117;
            end if;
        when multiplication_with_reduction_117 => 
            next_state <= multiplication_with_reduction_117;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_118;
            end if;
        when multiplication_with_reduction_118 => 
            next_state <= multiplication_with_reduction_118;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_119;
            end if;
        when multiplication_with_reduction_119 => 
            next_state <= multiplication_with_reduction_119;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_120;
            end if;
        when multiplication_with_reduction_120 => 
            next_state <= multiplication_with_reduction_120;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_121;
            end if;
        when multiplication_with_reduction_121 => 
            next_state <= multiplication_with_reduction_121;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_122;
            end if;
        when multiplication_with_reduction_122 => 
            next_state <= multiplication_with_reduction_122;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_123;
            end if;
        when multiplication_with_reduction_123 => 
            next_state <= multiplication_with_reduction_123;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_124;
            end if;
        when multiplication_with_reduction_124 => 
            next_state <= multiplication_with_reduction_124;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_125;
            end if;
        when multiplication_with_reduction_125 => 
            next_state <= multiplication_with_reduction_125;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_126;
            end if;
        when multiplication_with_reduction_126 => 
            next_state <= multiplication_with_reduction_126;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_127;
            end if;
        when multiplication_with_reduction_127 => 
            next_state <= multiplication_with_reduction_127;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_128;
            end if;
        when multiplication_with_reduction_128 => 
            next_state <= multiplication_with_reduction_128;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_129;
            end if;
        when multiplication_with_reduction_129 => 
            next_state <= multiplication_with_reduction_129;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_130;
            end if;
        when multiplication_with_reduction_130 => 
            next_state <= multiplication_with_reduction_130;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_131;
            end if;
        when multiplication_with_reduction_131 => 
            next_state <= multiplication_with_reduction_131;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_132;
            end if;
        when multiplication_with_reduction_132 => 
            next_state <= multiplication_with_reduction_132;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_133;
            end if;
        when multiplication_with_reduction_133 => 
            next_state <= multiplication_with_reduction_133;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_134;
            end if;
        when multiplication_with_reduction_134 => 
            next_state <= multiplication_with_reduction_134;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_135;
            end if;
        when multiplication_with_reduction_135 => 
            next_state <= multiplication_with_reduction_135;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_136;
            end if;
        when multiplication_with_reduction_136 => 
            next_state <= multiplication_with_reduction_136;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_137;
            end if;
        when multiplication_with_reduction_137 => 
            next_state <= multiplication_with_reduction_137;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_138;
            end if;
        when multiplication_with_reduction_138 => 
            next_state <= multiplication_with_reduction_138;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_139;
            end if;
        when multiplication_with_reduction_139 => 
            next_state <= multiplication_with_reduction_139;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_140;
            end if;
        when multiplication_with_reduction_140 => 
            next_state <= multiplication_with_reduction_140;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_141;
            end if;
        when multiplication_with_reduction_141 => 
            next_state <= multiplication_with_reduction_141;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_142;
            end if;
        when multiplication_with_reduction_142 => 
            next_state <= multiplication_with_reduction_142;
            if(ultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when multiplication_with_reduction_144 => 
            next_state <= multiplication_with_reduction_144;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_145;
            end if;
        when multiplication_with_reduction_145 => 
            next_state <= multiplication_with_reduction_145;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_146;
            end if;
        when multiplication_with_reduction_146 => 
            next_state <= multiplication_with_reduction_146;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_147;
            end if;
        when multiplication_with_reduction_147 => 
            next_state <= multiplication_with_reduction_147;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_148;
            end if;
        when multiplication_with_reduction_148 => 
            next_state <= multiplication_with_reduction_148;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_149;
            end if;
        when multiplication_with_reduction_149 => 
            next_state <= multiplication_with_reduction_149;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_150;
            end if;
        when multiplication_with_reduction_150 => 
            next_state <= multiplication_with_reduction_150;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_151;
            end if;
        when multiplication_with_reduction_151 => 
            next_state <= multiplication_with_reduction_151;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_152;
            end if;
        when multiplication_with_reduction_152 => 
            next_state <= multiplication_with_reduction_152;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_153;
            end if;
        when multiplication_with_reduction_153 => 
            next_state <= multiplication_with_reduction_153;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_154;
            end if;
        when multiplication_with_reduction_154 => 
            next_state <= multiplication_with_reduction_154;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_155;
            end if;
        when multiplication_with_reduction_155 => 
            next_state <= multiplication_with_reduction_155;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_156;
            end if;
        when multiplication_with_reduction_156 => 
            next_state <= multiplication_with_reduction_156;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_157;
            end if;
        when multiplication_with_reduction_157 => 
            next_state <= multiplication_with_reduction_157;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_158;
            end if;
        when multiplication_with_reduction_158 => 
            next_state <= multiplication_with_reduction_158;
            if(ultimate_operation = '1') then
                if(operands_size = "110") then
                    next_state <= multiplication_with_reduction_159;
                else
                    next_state <= multiplication_with_reduction_206;
                end if;
            end if;
        when multiplication_with_reduction_159 => 
            next_state <= multiplication_with_reduction_159;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_160;
            end if;
        when multiplication_with_reduction_160 => 
            next_state <= multiplication_with_reduction_160;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_161;
            end if;
        when multiplication_with_reduction_161 => 
            next_state <= multiplication_with_reduction_161;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_162;
            end if;
        when multiplication_with_reduction_162 => 
            next_state <= multiplication_with_reduction_162;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_163;
            end if;
        when multiplication_with_reduction_163 => 
            next_state <= multiplication_with_reduction_163;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_164;
            end if;
        when multiplication_with_reduction_164 => 
            next_state <= multiplication_with_reduction_164;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_165;
            end if;
        when multiplication_with_reduction_165 => 
            next_state <= multiplication_with_reduction_165;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_166;
            end if;
        when multiplication_with_reduction_166 => 
            next_state <= multiplication_with_reduction_166;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_167;
            end if;
        when multiplication_with_reduction_167 => 
            next_state <= multiplication_with_reduction_167;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_168;
            end if;
        when multiplication_with_reduction_168 => 
            next_state <= multiplication_with_reduction_168;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_169;
            end if;
        when multiplication_with_reduction_169 => 
            next_state <= multiplication_with_reduction_169;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_170;
            end if;
        when multiplication_with_reduction_170 => 
            next_state <= multiplication_with_reduction_170;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_171;
            end if;
        when multiplication_with_reduction_171 => 
            next_state <= multiplication_with_reduction_171;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_172;
            end if;
        when multiplication_with_reduction_172 => 
            next_state <= multiplication_with_reduction_172;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_173;
            end if;
        when multiplication_with_reduction_173 => 
            next_state <= multiplication_with_reduction_173;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_174;
            end if;
        when multiplication_with_reduction_174 => 
            next_state <= multiplication_with_reduction_174;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_175;
            end if;
        when multiplication_with_reduction_175 => 
            next_state <= multiplication_with_reduction_175;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_176;
            end if;
        when multiplication_with_reduction_176 => 
            next_state <= multiplication_with_reduction_176;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_177;
            end if;
        when multiplication_with_reduction_177 => 
            next_state <= multiplication_with_reduction_177;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_178;
            end if;
        when multiplication_with_reduction_178 => 
            next_state <= multiplication_with_reduction_178;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_179;
            end if;
        when multiplication_with_reduction_179 => 
            next_state <= multiplication_with_reduction_179;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_180;
            end if;
        when multiplication_with_reduction_180 => 
            next_state <= multiplication_with_reduction_180;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_181;
            end if;
        when multiplication_with_reduction_181 => 
            next_state <= multiplication_with_reduction_181;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_182;
            end if;
        when multiplication_with_reduction_182 => 
            next_state <= multiplication_with_reduction_182;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_183;
            end if;
        when multiplication_with_reduction_183 => 
            next_state <= multiplication_with_reduction_183;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_184;
            end if;
        when multiplication_with_reduction_184 => 
            next_state <= multiplication_with_reduction_184;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_185;
            end if;
        when multiplication_with_reduction_185 => 
            next_state <= multiplication_with_reduction_185;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_186;
            end if;
        when multiplication_with_reduction_186 => 
            next_state <= multiplication_with_reduction_186;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_187;
            end if;
        when multiplication_with_reduction_187 => 
            next_state <= multiplication_with_reduction_187;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_188;
            end if;
        when multiplication_with_reduction_188 => 
            next_state <= multiplication_with_reduction_188;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_189;
            end if;
        when multiplication_with_reduction_189 => 
            next_state <= multiplication_with_reduction_189;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_190;
            end if;
        when multiplication_with_reduction_190 => 
            next_state <= multiplication_with_reduction_190;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_191;
            end if;
        when multiplication_with_reduction_191 => 
            next_state <= multiplication_with_reduction_191;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_192;
            end if;
        when multiplication_with_reduction_192 => 
            next_state <= multiplication_with_reduction_192;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_193;
            end if;
        when multiplication_with_reduction_193 => 
            next_state <= multiplication_with_reduction_193;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_194;
            end if;
        when multiplication_with_reduction_194 => 
            next_state <= multiplication_with_reduction_194;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_195;
            end if;
        when multiplication_with_reduction_195 => 
            next_state <= multiplication_with_reduction_195;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_196;
            end if;
        when multiplication_with_reduction_196 => 
            next_state <= multiplication_with_reduction_196;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_197;
            end if;
        when multiplication_with_reduction_197 => 
            next_state <= multiplication_with_reduction_197;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_198;
            end if;
        when multiplication_with_reduction_198 => 
            next_state <= multiplication_with_reduction_198;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_199;
            end if;
        when multiplication_with_reduction_199 => 
            next_state <= multiplication_with_reduction_199;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_200;
            end if;
        when multiplication_with_reduction_200 => 
            next_state <= multiplication_with_reduction_200;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_201;
            end if;
        when multiplication_with_reduction_201 => 
            next_state <= multiplication_with_reduction_201;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_202;
            end if;
        when multiplication_with_reduction_202 => 
            next_state <= multiplication_with_reduction_202;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_203;
            end if;
        when multiplication_with_reduction_203 => 
            next_state <= multiplication_with_reduction_203;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_204;
            end if;
        when multiplication_with_reduction_204 => 
            next_state <= multiplication_with_reduction_204;
            if(ultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when multiplication_with_reduction_206 => 
            next_state <= multiplication_with_reduction_206;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_207;
            end if;
        when multiplication_with_reduction_207 => 
            next_state <= multiplication_with_reduction_207;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_208;
            end if;
        when multiplication_with_reduction_208 => 
            next_state <= multiplication_with_reduction_208;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_209;
            end if;
        when multiplication_with_reduction_209 => 
            next_state <= multiplication_with_reduction_209;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_210;
            end if;
        when multiplication_with_reduction_210 => 
            next_state <= multiplication_with_reduction_210;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_211;
            end if;
        when multiplication_with_reduction_211 => 
            next_state <= multiplication_with_reduction_211;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_212;
            end if;
        when multiplication_with_reduction_212 => 
            next_state <= multiplication_with_reduction_212;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_213;
            end if;
        when multiplication_with_reduction_213 => 
            next_state <= multiplication_with_reduction_213;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_214;
            end if;
        when multiplication_with_reduction_214 => 
            next_state <= multiplication_with_reduction_214;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_215;
            end if;
        when multiplication_with_reduction_215 => 
            next_state <= multiplication_with_reduction_215;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_216;
            end if;
        when multiplication_with_reduction_216 => 
            next_state <= multiplication_with_reduction_216;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_217;
            end if;
        when multiplication_with_reduction_217 => 
            next_state <= multiplication_with_reduction_217;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_218;
            end if;
        when multiplication_with_reduction_218 => 
            next_state <= multiplication_with_reduction_218;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_219;
            end if;
        when multiplication_with_reduction_219 => 
            next_state <= multiplication_with_reduction_219;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_220;
            end if;
        when multiplication_with_reduction_220 => 
            next_state <= multiplication_with_reduction_220;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_221;
            end if;
        when multiplication_with_reduction_221 => 
            next_state <= multiplication_with_reduction_221;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_222;
            end if;
        when multiplication_with_reduction_222 => 
            next_state <= multiplication_with_reduction_222;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_223;
            end if;
        when multiplication_with_reduction_223 => 
            next_state <= multiplication_with_reduction_223;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_224;
            end if;
        when multiplication_with_reduction_224 => 
            next_state <= multiplication_with_reduction_224;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_225;
            end if;
        when multiplication_with_reduction_225 => 
            next_state <= multiplication_with_reduction_225;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_226;
            end if;
        when multiplication_with_reduction_226 => 
            next_state <= multiplication_with_reduction_226;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_227;
            end if;
        when multiplication_with_reduction_227 => 
            next_state <= multiplication_with_reduction_227;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_228;
            end if;
        when multiplication_with_reduction_228 => 
            next_state <= multiplication_with_reduction_228;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_229;
            end if;
        when multiplication_with_reduction_229 => 
            next_state <= multiplication_with_reduction_229;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_230;
            end if;
        when multiplication_with_reduction_230 => 
            next_state <= multiplication_with_reduction_230;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_231;
            end if;
        when multiplication_with_reduction_231 => 
            next_state <= multiplication_with_reduction_231;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_232;
            end if;
        when multiplication_with_reduction_232 => 
            next_state <= multiplication_with_reduction_232;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_233;
            end if;
        when multiplication_with_reduction_233 => 
            next_state <= multiplication_with_reduction_233;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_234;
            end if;
        when multiplication_with_reduction_234 => 
            next_state <= multiplication_with_reduction_234;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_235;
            end if;
        when multiplication_with_reduction_235 => 
            next_state <= multiplication_with_reduction_235;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_236;
            end if;
        when multiplication_with_reduction_236 => 
            next_state <= multiplication_with_reduction_236;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_237;
            end if;
        when multiplication_with_reduction_237 => 
            next_state <= multiplication_with_reduction_237;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_238;
            end if;
        when multiplication_with_reduction_238 => 
            next_state <= multiplication_with_reduction_238;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_239;
            end if;
        when multiplication_with_reduction_239 => 
            next_state <= multiplication_with_reduction_239;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_240;
            end if;
        when multiplication_with_reduction_240 => 
            next_state <= multiplication_with_reduction_240;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_241;
            end if;
        when multiplication_with_reduction_241 => 
            next_state <= multiplication_with_reduction_241;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_242;
            end if;
        when multiplication_with_reduction_242 => 
            next_state <= multiplication_with_reduction_242;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_243;
            end if;
        when multiplication_with_reduction_243 => 
            next_state <= multiplication_with_reduction_243;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_244;
            end if;
        when multiplication_with_reduction_244 => 
            next_state <= multiplication_with_reduction_244;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_245;
            end if;
        when multiplication_with_reduction_245 => 
            next_state <= multiplication_with_reduction_245;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_246;
            end if;
        when multiplication_with_reduction_246 => 
            next_state <= multiplication_with_reduction_246;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_247;
            end if;
        when multiplication_with_reduction_247 => 
            next_state <= multiplication_with_reduction_247;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_248;
            end if;
        when multiplication_with_reduction_248 => 
            next_state <= multiplication_with_reduction_248;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_249;
            end if;
        when multiplication_with_reduction_249 => 
            next_state <= multiplication_with_reduction_249;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_250;
            end if;
        when multiplication_with_reduction_250 => 
            next_state <= multiplication_with_reduction_250;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_251;
            end if;
        when multiplication_with_reduction_251 => 
            next_state <= multiplication_with_reduction_251;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_252;
            end if;
        when multiplication_with_reduction_252 => 
            next_state <= multiplication_with_reduction_252;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_253;
            end if;
        when multiplication_with_reduction_253 => 
            next_state <= multiplication_with_reduction_253;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_254;
            end if;
        when multiplication_with_reduction_254 => 
            next_state <= multiplication_with_reduction_254;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_255;
            end if;
        when multiplication_with_reduction_255 => 
            next_state <= multiplication_with_reduction_255;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_256;
            end if;
        when multiplication_with_reduction_256 => 
            next_state <= multiplication_with_reduction_256;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_257;
            end if;
        when multiplication_with_reduction_257 => 
            next_state <= multiplication_with_reduction_257;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_258;
            end if;
        when multiplication_with_reduction_258 => 
            next_state <= multiplication_with_reduction_258;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_259;
            end if;
        when multiplication_with_reduction_259 => 
            next_state <= multiplication_with_reduction_259;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_260;
            end if;
        when multiplication_with_reduction_260 => 
            next_state <= multiplication_with_reduction_260;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_261;
            end if;
        when multiplication_with_reduction_261 => 
            next_state <= multiplication_with_reduction_261;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_262;
            end if;
        when multiplication_with_reduction_262 => 
            next_state <= multiplication_with_reduction_262;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_263;
            end if;
        when multiplication_with_reduction_263 => 
            next_state <= multiplication_with_reduction_263;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_264;
            end if;
        when multiplication_with_reduction_264 => 
            next_state <= multiplication_with_reduction_264;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_265;
            end if;
        when multiplication_with_reduction_265 => 
            next_state <= multiplication_with_reduction_265;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_266;
            end if;
        when multiplication_with_reduction_266 => 
            next_state <= multiplication_with_reduction_266;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_267;
            end if;
        when multiplication_with_reduction_267 => 
            next_state <= multiplication_with_reduction_267;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_268;
            end if;
        when multiplication_with_reduction_268 => 
            next_state <= multiplication_with_reduction_268;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_269;
            end if;
        when multiplication_with_reduction_269 => 
            next_state <= multiplication_with_reduction_269;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_270;
            end if;
        when multiplication_with_reduction_270 => 
            next_state <= multiplication_with_reduction_270;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_271;
            end if;
        when multiplication_with_reduction_271 => 
            next_state <= multiplication_with_reduction_271;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_272;
            end if;
        when multiplication_with_reduction_272 => 
            next_state <= multiplication_with_reduction_272;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_273;
            end if;
        when multiplication_with_reduction_273 => 
            next_state <= multiplication_with_reduction_273;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_274;
            end if;
        when multiplication_with_reduction_274 => 
            next_state <= multiplication_with_reduction_274;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_275;
            end if;
        when multiplication_with_reduction_275 => 
            next_state <= multiplication_with_reduction_275;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_276;
            end if;
        when multiplication_with_reduction_276 => 
            next_state <= multiplication_with_reduction_276;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_277;
            end if;
        when multiplication_with_reduction_277 => 
            next_state <= multiplication_with_reduction_277;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_278;
            end if;
        when multiplication_with_reduction_278 => 
            next_state <= multiplication_with_reduction_278;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_279;
            end if;
        when multiplication_with_reduction_279 => 
            next_state <= multiplication_with_reduction_279;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_280;
            end if;
        when multiplication_with_reduction_280 => 
            next_state <= multiplication_with_reduction_280;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_281;
            end if;
        when multiplication_with_reduction_281 => 
            next_state <= multiplication_with_reduction_281;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_282;
            end if;
        when multiplication_with_reduction_282 => 
            next_state <= multiplication_with_reduction_282;
            if(ultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when multiplication_with_reduction_special_prime_1_0 => 
            next_state <= multiplication_with_reduction_special_prime_1_0;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_1;
            end if;
        when multiplication_with_reduction_special_prime_1_1 => 
            next_state <= multiplication_with_reduction_special_prime_1_1;
            if(ultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when multiplication_with_reduction_special_prime_1_3 => 
            next_state <= multiplication_with_reduction_special_prime_1_3;
            if(ultimate_operation = '1') then
                if(operands_size = "001") then
                    next_state <= multiplication_with_reduction_special_prime_1_4;
                else
                    next_state <= multiplication_with_reduction_special_prime_1_10;
                end if;
            end if;
        when multiplication_with_reduction_special_prime_1_4 => 
            next_state <= multiplication_with_reduction_special_prime_1_4;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_5;
            end if;
        when multiplication_with_reduction_special_prime_1_5 => 
            next_state <= multiplication_with_reduction_special_prime_1_5;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_6;
            end if;
        when multiplication_with_reduction_special_prime_1_6 => 
            next_state <= multiplication_with_reduction_special_prime_1_6;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_7;
            end if;
        when multiplication_with_reduction_special_prime_1_7 => 
            next_state <= multiplication_with_reduction_special_prime_1_7;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_8;
            end if;
        when multiplication_with_reduction_special_prime_1_8 => 
            next_state <= multiplication_with_reduction_special_prime_1_8;
            if(ultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when multiplication_with_reduction_special_prime_1_10 => 
            next_state <= multiplication_with_reduction_special_prime_1_10;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_11;
            end if;
        when multiplication_with_reduction_special_prime_1_11 => 
            next_state <= multiplication_with_reduction_special_prime_1_11;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_12;
            end if;
        when multiplication_with_reduction_special_prime_1_12 => 
            next_state <= multiplication_with_reduction_special_prime_1_12;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_13;
            end if;
        when multiplication_with_reduction_special_prime_1_13 => 
            next_state <= multiplication_with_reduction_special_prime_1_13;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_14;
            end if;
        when multiplication_with_reduction_special_prime_1_14 => 
            next_state <= multiplication_with_reduction_special_prime_1_14;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_15;
            end if;
        when multiplication_with_reduction_special_prime_1_15 => 
            next_state <= multiplication_with_reduction_special_prime_1_15;
            if(ultimate_operation = '1') then
                if(operands_size = "010") then
                    next_state <= multiplication_with_reduction_special_prime_1_16;
                else
                    next_state <= multiplication_with_reduction_special_prime_1_25;
                end if;
            end if;
        when multiplication_with_reduction_special_prime_1_16 => 
            next_state <= multiplication_with_reduction_special_prime_1_16;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_17;
            end if;
        when multiplication_with_reduction_special_prime_1_17 => 
            next_state <= multiplication_with_reduction_special_prime_1_17;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_18;
            end if;
        when multiplication_with_reduction_special_prime_1_18 => 
            next_state <= multiplication_with_reduction_special_prime_1_18;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_19;
            end if;
        when multiplication_with_reduction_special_prime_1_19 => 
            next_state <= multiplication_with_reduction_special_prime_1_19;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_20;
            end if;
        when multiplication_with_reduction_special_prime_1_20 => 
            next_state <= multiplication_with_reduction_special_prime_1_20;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_21;
            end if;
        when multiplication_with_reduction_special_prime_1_21 => 
            next_state <= multiplication_with_reduction_special_prime_1_21;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_22;
            end if;
        when multiplication_with_reduction_special_prime_1_22 => 
            next_state <= multiplication_with_reduction_special_prime_1_22;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_23;
            end if;
        when multiplication_with_reduction_special_prime_1_23 => 
            next_state <= multiplication_with_reduction_special_prime_1_23;
            if(ultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when multiplication_with_reduction_special_prime_1_25 => 
            next_state <= multiplication_with_reduction_special_prime_1_25;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_26;
            end if;
        when multiplication_with_reduction_special_prime_1_26 => 
            next_state <= multiplication_with_reduction_special_prime_1_26;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_27;
            end if;
        when multiplication_with_reduction_special_prime_1_27 => 
            next_state <= multiplication_with_reduction_special_prime_1_27;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_28;
            end if;
        when multiplication_with_reduction_special_prime_1_28 => 
            next_state <= multiplication_with_reduction_special_prime_1_28;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_29;
            end if;
        when multiplication_with_reduction_special_prime_1_29 => 
            next_state <= multiplication_with_reduction_special_prime_1_29;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_30;
            end if;
        when multiplication_with_reduction_special_prime_1_30 => 
            next_state <= multiplication_with_reduction_special_prime_1_30;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_31;
            end if;
        when multiplication_with_reduction_special_prime_1_31 => 
            next_state <= multiplication_with_reduction_special_prime_1_31;
            if(ultimate_operation = '1') then
                if(operands_size = "011") then
                    next_state <= multiplication_with_reduction_special_prime_1_32;
                else
                    next_state <= multiplication_with_reduction_special_prime_1_47;
                end if;
            end if;
        when multiplication_with_reduction_special_prime_1_32 => 
            next_state <= multiplication_with_reduction_special_prime_1_32;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_33;
            end if;
        when multiplication_with_reduction_special_prime_1_33 => 
            next_state <= multiplication_with_reduction_special_prime_1_33;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_34;
            end if;
        when multiplication_with_reduction_special_prime_1_34 => 
            next_state <= multiplication_with_reduction_special_prime_1_34;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_35;
            end if;
        when multiplication_with_reduction_special_prime_1_35 => 
            next_state <= multiplication_with_reduction_special_prime_1_35;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_36;
            end if;
        when multiplication_with_reduction_special_prime_1_36 => 
            next_state <= multiplication_with_reduction_special_prime_1_36;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_37;
            end if;
        when multiplication_with_reduction_special_prime_1_37 => 
            next_state <= multiplication_with_reduction_special_prime_1_37;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_38;
            end if;
        when multiplication_with_reduction_special_prime_1_38 => 
            next_state <= multiplication_with_reduction_special_prime_1_38;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_39;
            end if;
        when multiplication_with_reduction_special_prime_1_39 => 
            next_state <= multiplication_with_reduction_special_prime_1_39;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_40;
            end if;
        when multiplication_with_reduction_special_prime_1_40 => 
            next_state <= multiplication_with_reduction_special_prime_1_40;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_41;
            end if;
        when multiplication_with_reduction_special_prime_1_41 => 
            next_state <= multiplication_with_reduction_special_prime_1_41;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_42;
            end if;
        when multiplication_with_reduction_special_prime_1_42 => 
            next_state <= multiplication_with_reduction_special_prime_1_42;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_43;
            end if;
        when multiplication_with_reduction_special_prime_1_43 => 
            next_state <= multiplication_with_reduction_special_prime_1_43;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_44;
            end if;
        when multiplication_with_reduction_special_prime_1_44 => 
            next_state <= multiplication_with_reduction_special_prime_1_44;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_45;
            end if;
        when multiplication_with_reduction_special_prime_1_45 => 
            next_state <= multiplication_with_reduction_special_prime_1_45;
            if(ultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when multiplication_with_reduction_special_prime_1_47 =>
            next_state <= multiplication_with_reduction_special_prime_1_47;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_48;
            end if;
        when multiplication_with_reduction_special_prime_1_48 =>
            next_state <= multiplication_with_reduction_special_prime_1_48;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_49;
            end if;
        when multiplication_with_reduction_special_prime_1_49 =>
            next_state <= multiplication_with_reduction_special_prime_1_49;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_50;
            end if;
        when multiplication_with_reduction_special_prime_1_50 =>
            next_state <= multiplication_with_reduction_special_prime_1_50;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_51;
            end if;
        when multiplication_with_reduction_special_prime_1_51 =>
            next_state <= multiplication_with_reduction_special_prime_1_51;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_52;
            end if;
        when multiplication_with_reduction_special_prime_1_52 =>
            next_state <= multiplication_with_reduction_special_prime_1_52;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_53;
            end if;
        when multiplication_with_reduction_special_prime_1_53 =>
            next_state <= multiplication_with_reduction_special_prime_1_53;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_54;
            end if;
        when multiplication_with_reduction_special_prime_1_54 =>
            next_state <= multiplication_with_reduction_special_prime_1_54;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_55;
            end if;
        when multiplication_with_reduction_special_prime_1_55 =>
            next_state <= multiplication_with_reduction_special_prime_1_55;
            if(ultimate_operation = '1') then
                if(operands_size = "100") then
                    next_state <= multiplication_with_reduction_special_prime_1_56;
                else
                    next_state <= multiplication_with_reduction_special_prime_1_79;
                end if;
            end if;
        when multiplication_with_reduction_special_prime_1_56 =>
            next_state <= multiplication_with_reduction_special_prime_1_56;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_57;
            end if;
        when multiplication_with_reduction_special_prime_1_57 =>
            next_state <= multiplication_with_reduction_special_prime_1_57;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_58;
            end if;
        when multiplication_with_reduction_special_prime_1_58 =>
            next_state <= multiplication_with_reduction_special_prime_1_58;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_59;
            end if;
        when multiplication_with_reduction_special_prime_1_59 =>
            next_state <= multiplication_with_reduction_special_prime_1_59;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_60;
            end if;
        when multiplication_with_reduction_special_prime_1_60 =>
            next_state <= multiplication_with_reduction_special_prime_1_60;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_61;
            end if;
        when multiplication_with_reduction_special_prime_1_61 =>
            next_state <= multiplication_with_reduction_special_prime_1_61;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_62;
            end if;
        when multiplication_with_reduction_special_prime_1_62 =>
            next_state <= multiplication_with_reduction_special_prime_1_62;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_63;
            end if;
        when multiplication_with_reduction_special_prime_1_63 =>
            next_state <= multiplication_with_reduction_special_prime_1_63;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_64;
            end if;
        when multiplication_with_reduction_special_prime_1_64 =>
            next_state <= multiplication_with_reduction_special_prime_1_64;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_65;
            end if;
        when multiplication_with_reduction_special_prime_1_65 =>
            next_state <= multiplication_with_reduction_special_prime_1_65;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_66;
            end if;
        when multiplication_with_reduction_special_prime_1_66 =>
            next_state <= multiplication_with_reduction_special_prime_1_66;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_67;
            end if;
        when multiplication_with_reduction_special_prime_1_67 =>
            next_state <= multiplication_with_reduction_special_prime_1_67;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_68;
            end if;
        when multiplication_with_reduction_special_prime_1_68 =>
            next_state <= multiplication_with_reduction_special_prime_1_68;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_69;
            end if;
        when multiplication_with_reduction_special_prime_1_69 =>
            next_state <= multiplication_with_reduction_special_prime_1_69;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_70;
            end if;
        when multiplication_with_reduction_special_prime_1_70 =>
            next_state <= multiplication_with_reduction_special_prime_1_70;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_71;
            end if;
        when multiplication_with_reduction_special_prime_1_71 =>
            next_state <= multiplication_with_reduction_special_prime_1_71;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_72;
            end if;
        when multiplication_with_reduction_special_prime_1_72 =>
            next_state <= multiplication_with_reduction_special_prime_1_72;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_73;
            end if;
        when multiplication_with_reduction_special_prime_1_73 =>
            next_state <= multiplication_with_reduction_special_prime_1_73;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_74;
            end if;
        when multiplication_with_reduction_special_prime_1_74 =>
            next_state <= multiplication_with_reduction_special_prime_1_74;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_75;
            end if;
        when multiplication_with_reduction_special_prime_1_75 =>
            next_state <= multiplication_with_reduction_special_prime_1_75;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_76;
            end if;
        when multiplication_with_reduction_special_prime_1_76 =>
            next_state <= multiplication_with_reduction_special_prime_1_76;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_77;
            end if;
        when multiplication_with_reduction_special_prime_1_77 =>
            next_state <= multiplication_with_reduction_special_prime_1_77;
            if(ultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when multiplication_with_reduction_special_prime_1_79 =>
            next_state <= multiplication_with_reduction_special_prime_1_79;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_80;
            end if;
        when multiplication_with_reduction_special_prime_1_80 =>
            next_state <= multiplication_with_reduction_special_prime_1_80;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_81;
            end if;
        when multiplication_with_reduction_special_prime_1_81 =>
            next_state <= multiplication_with_reduction_special_prime_1_81;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_82;
            end if;
        when multiplication_with_reduction_special_prime_1_82 =>
            next_state <= multiplication_with_reduction_special_prime_1_82;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_83;
            end if;
        when multiplication_with_reduction_special_prime_1_83 =>
            next_state <= multiplication_with_reduction_special_prime_1_83;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_84;
            end if;
        when multiplication_with_reduction_special_prime_1_84 =>
            next_state <= multiplication_with_reduction_special_prime_1_84;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_85;
            end if;
        when multiplication_with_reduction_special_prime_1_85 =>
            next_state <= multiplication_with_reduction_special_prime_1_85;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_86;
            end if;
        when multiplication_with_reduction_special_prime_1_86 =>
            next_state <= multiplication_with_reduction_special_prime_1_86;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_87;
            end if;
        when multiplication_with_reduction_special_prime_1_87 =>
            next_state <= multiplication_with_reduction_special_prime_1_87;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_88;
            end if;
        when multiplication_with_reduction_special_prime_1_88 =>
            next_state <= multiplication_with_reduction_special_prime_1_88;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_89;
            end if;
        when multiplication_with_reduction_special_prime_1_89 =>
            next_state <= multiplication_with_reduction_special_prime_1_89;
            if(ultimate_operation = '1') then
                if(operands_size = "101") then
                    next_state <= multiplication_with_reduction_special_prime_1_90;
                else
                    next_state <= multiplication_with_reduction_special_prime_1_123;
                end if;
            end if;
        when multiplication_with_reduction_special_prime_1_90 =>
            next_state <= multiplication_with_reduction_special_prime_1_90;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_91;
            end if;
        when multiplication_with_reduction_special_prime_1_91 =>
            next_state <= multiplication_with_reduction_special_prime_1_91;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_92;
            end if;
        when multiplication_with_reduction_special_prime_1_92 =>
            next_state <= multiplication_with_reduction_special_prime_1_92;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_93;
            end if;
        when multiplication_with_reduction_special_prime_1_93 =>
            next_state <= multiplication_with_reduction_special_prime_1_93;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_94;
            end if;
        when multiplication_with_reduction_special_prime_1_94 =>
            next_state <= multiplication_with_reduction_special_prime_1_94;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_95;
            end if;
        when multiplication_with_reduction_special_prime_1_95 =>
            next_state <= multiplication_with_reduction_special_prime_1_95;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_96;
            end if;
        when multiplication_with_reduction_special_prime_1_96 =>
            next_state <= multiplication_with_reduction_special_prime_1_96;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_97;
            end if;
        when multiplication_with_reduction_special_prime_1_97 =>
            next_state <= multiplication_with_reduction_special_prime_1_97;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_98;
            end if;
        when multiplication_with_reduction_special_prime_1_98 =>
            next_state <= multiplication_with_reduction_special_prime_1_98;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_99;
            end if;
        when multiplication_with_reduction_special_prime_1_99 =>
            next_state <= multiplication_with_reduction_special_prime_1_99;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_100;
            end if;
        when multiplication_with_reduction_special_prime_1_100 =>
            next_state <= multiplication_with_reduction_special_prime_1_100;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_101;
            end if;
        when multiplication_with_reduction_special_prime_1_101 =>
            next_state <= multiplication_with_reduction_special_prime_1_101;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_102;
            end if;
        when multiplication_with_reduction_special_prime_1_102 =>
            next_state <= multiplication_with_reduction_special_prime_1_102;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_103;
            end if;
        when multiplication_with_reduction_special_prime_1_103 =>
            next_state <= multiplication_with_reduction_special_prime_1_103;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_104;
            end if;
        when multiplication_with_reduction_special_prime_1_104 =>
            next_state <= multiplication_with_reduction_special_prime_1_104;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_105;
            end if;
        when multiplication_with_reduction_special_prime_1_105 =>
            next_state <= multiplication_with_reduction_special_prime_1_105;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_106;
            end if;
        when multiplication_with_reduction_special_prime_1_106 =>
            next_state <= multiplication_with_reduction_special_prime_1_106;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_107;
            end if;
        when multiplication_with_reduction_special_prime_1_107 =>
            next_state <= multiplication_with_reduction_special_prime_1_107;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_108;
            end if;
        when multiplication_with_reduction_special_prime_1_108 =>
            next_state <= multiplication_with_reduction_special_prime_1_108;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_109;
            end if;
        when multiplication_with_reduction_special_prime_1_109 =>
            next_state <= multiplication_with_reduction_special_prime_1_109;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_110;
            end if;
        when multiplication_with_reduction_special_prime_1_110 =>
            next_state <= multiplication_with_reduction_special_prime_1_110;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_111;
            end if;
        when multiplication_with_reduction_special_prime_1_111 =>
            next_state <= multiplication_with_reduction_special_prime_1_111;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_112;
            end if;
        when multiplication_with_reduction_special_prime_1_112 =>
            next_state <= multiplication_with_reduction_special_prime_1_112;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_113;
            end if;
        when multiplication_with_reduction_special_prime_1_113 =>
            next_state <= multiplication_with_reduction_special_prime_1_113;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_114;
            end if;
        when multiplication_with_reduction_special_prime_1_114 =>
            next_state <= multiplication_with_reduction_special_prime_1_114;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_115;
            end if;
        when multiplication_with_reduction_special_prime_1_115 =>
            next_state <= multiplication_with_reduction_special_prime_1_115;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_116;
            end if;
        when multiplication_with_reduction_special_prime_1_116 =>
            next_state <= multiplication_with_reduction_special_prime_1_116;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_117;
            end if;
        when multiplication_with_reduction_special_prime_1_117 =>
            next_state <= multiplication_with_reduction_special_prime_1_117;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_118;
            end if;
        when multiplication_with_reduction_special_prime_1_118 =>
            next_state <= multiplication_with_reduction_special_prime_1_118;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_119;
            end if;
        when multiplication_with_reduction_special_prime_1_119 =>
            next_state <= multiplication_with_reduction_special_prime_1_119;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_120;
            end if;
        when multiplication_with_reduction_special_prime_1_120 =>
            next_state <= multiplication_with_reduction_special_prime_1_120;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_121;
            end if;
        when multiplication_with_reduction_special_prime_1_121 =>
            next_state <= multiplication_with_reduction_special_prime_1_121;
            if(ultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when multiplication_with_reduction_special_prime_1_123 =>
            next_state <= multiplication_with_reduction_special_prime_1_123;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_124;
            end if;
        when multiplication_with_reduction_special_prime_1_124 =>
            next_state <= multiplication_with_reduction_special_prime_1_124;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_125;
            end if;
        when multiplication_with_reduction_special_prime_1_125 =>
            next_state <= multiplication_with_reduction_special_prime_1_125;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_126;
            end if;
        when multiplication_with_reduction_special_prime_1_126 =>
            next_state <= multiplication_with_reduction_special_prime_1_126;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_127;
            end if;
        when multiplication_with_reduction_special_prime_1_127 =>
            next_state <= multiplication_with_reduction_special_prime_1_127;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_128;
            end if;
        when multiplication_with_reduction_special_prime_1_128 =>
            next_state <= multiplication_with_reduction_special_prime_1_128;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_129;
            end if;
        when multiplication_with_reduction_special_prime_1_129 =>
            next_state <= multiplication_with_reduction_special_prime_1_129;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_130;
            end if;
        when multiplication_with_reduction_special_prime_1_130 =>
            next_state <= multiplication_with_reduction_special_prime_1_130;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_131;
            end if;
        when multiplication_with_reduction_special_prime_1_131 =>
            next_state <= multiplication_with_reduction_special_prime_1_131;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_132;
            end if;
        when multiplication_with_reduction_special_prime_1_132 =>
            next_state <= multiplication_with_reduction_special_prime_1_132;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_133;
            end if;
        when multiplication_with_reduction_special_prime_1_133 =>
            next_state <= multiplication_with_reduction_special_prime_1_133;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_134;
            end if;
        when multiplication_with_reduction_special_prime_1_134 =>
            next_state <= multiplication_with_reduction_special_prime_1_134;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_135;
            end if;
        when multiplication_with_reduction_special_prime_1_135 =>
            next_state <= multiplication_with_reduction_special_prime_1_135;
            if(ultimate_operation = '1') then
                if(operands_size = "110")then
                    next_state <= multiplication_with_reduction_special_prime_1_136;
                else
                    next_state <= multiplication_with_reduction_special_prime_1_181;
                end if;
            end if;
        when multiplication_with_reduction_special_prime_1_136 =>
            next_state <= multiplication_with_reduction_special_prime_1_136;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_137;
            end if;
        when multiplication_with_reduction_special_prime_1_137 =>
            next_state <= multiplication_with_reduction_special_prime_1_137;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_138;
            end if;
        when multiplication_with_reduction_special_prime_1_138 =>
            next_state <= multiplication_with_reduction_special_prime_1_138;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_139;
            end if;
        when multiplication_with_reduction_special_prime_1_139 =>
            next_state <= multiplication_with_reduction_special_prime_1_139;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_140;
            end if;
        when multiplication_with_reduction_special_prime_1_140 =>
            next_state <= multiplication_with_reduction_special_prime_1_140;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_141;
            end if;
        when multiplication_with_reduction_special_prime_1_141 =>
            next_state <= multiplication_with_reduction_special_prime_1_141;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_142;
            end if;
        when multiplication_with_reduction_special_prime_1_142 =>
            next_state <= multiplication_with_reduction_special_prime_1_142;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_143;
            end if;
        when multiplication_with_reduction_special_prime_1_143 =>
            next_state <= multiplication_with_reduction_special_prime_1_143;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_144;
            end if;
        when multiplication_with_reduction_special_prime_1_144 =>
            next_state <= multiplication_with_reduction_special_prime_1_144;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_145;
            end if;
        when multiplication_with_reduction_special_prime_1_145 =>
            next_state <= multiplication_with_reduction_special_prime_1_145;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_146;
            end if;
        when multiplication_with_reduction_special_prime_1_146 =>
            next_state <= multiplication_with_reduction_special_prime_1_146;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_147;
            end if;
        when multiplication_with_reduction_special_prime_1_147 =>
            next_state <= multiplication_with_reduction_special_prime_1_147;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_148;
            end if;
        when multiplication_with_reduction_special_prime_1_148 =>
            next_state <= multiplication_with_reduction_special_prime_1_148;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_149;
            end if;
        when multiplication_with_reduction_special_prime_1_149 =>
            next_state <= multiplication_with_reduction_special_prime_1_149;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_150;
            end if;
        when multiplication_with_reduction_special_prime_1_150 =>
            next_state <= multiplication_with_reduction_special_prime_1_150;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_151;
            end if;
        when multiplication_with_reduction_special_prime_1_151 =>
            next_state <= multiplication_with_reduction_special_prime_1_151;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_152;
            end if;
        when multiplication_with_reduction_special_prime_1_152 =>
            next_state <= multiplication_with_reduction_special_prime_1_152;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_153;
            end if;
        when multiplication_with_reduction_special_prime_1_153 =>
            next_state <= multiplication_with_reduction_special_prime_1_153;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_154;
            end if;
        when multiplication_with_reduction_special_prime_1_154 =>
            next_state <= multiplication_with_reduction_special_prime_1_154;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_155;
            end if;
        when multiplication_with_reduction_special_prime_1_155 =>
            next_state <= multiplication_with_reduction_special_prime_1_155;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_156;
            end if;
        when multiplication_with_reduction_special_prime_1_156 =>
            next_state <= multiplication_with_reduction_special_prime_1_156;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_157;
            end if;
        when multiplication_with_reduction_special_prime_1_157 =>
            next_state <= multiplication_with_reduction_special_prime_1_157;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_158;
            end if;
        when multiplication_with_reduction_special_prime_1_158 =>
            next_state <= multiplication_with_reduction_special_prime_1_158;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_159;
            end if;
        when multiplication_with_reduction_special_prime_1_159 =>
            next_state <= multiplication_with_reduction_special_prime_1_159;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_160;
            end if;
        when multiplication_with_reduction_special_prime_1_160 =>
            next_state <= multiplication_with_reduction_special_prime_1_160;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_161;
            end if;
        when multiplication_with_reduction_special_prime_1_161 =>
            next_state <= multiplication_with_reduction_special_prime_1_161;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_162;
            end if;
        when multiplication_with_reduction_special_prime_1_162 =>
            next_state <= multiplication_with_reduction_special_prime_1_162;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_163;
            end if;
        when multiplication_with_reduction_special_prime_1_163 =>
            next_state <= multiplication_with_reduction_special_prime_1_163;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_164;
            end if;
        when multiplication_with_reduction_special_prime_1_164 =>
            next_state <= multiplication_with_reduction_special_prime_1_164;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_165;
            end if;
        when multiplication_with_reduction_special_prime_1_165 =>
            next_state <= multiplication_with_reduction_special_prime_1_165;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_166;
            end if;
        when multiplication_with_reduction_special_prime_1_166 =>
            next_state <= multiplication_with_reduction_special_prime_1_166;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_167;
            end if;
        when multiplication_with_reduction_special_prime_1_167 =>
            next_state <= multiplication_with_reduction_special_prime_1_167;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_168;
            end if;
        when multiplication_with_reduction_special_prime_1_168 =>
            next_state <= multiplication_with_reduction_special_prime_1_168;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_169;
            end if;
        when multiplication_with_reduction_special_prime_1_169 =>
            next_state <= multiplication_with_reduction_special_prime_1_169;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_170;
            end if;
        when multiplication_with_reduction_special_prime_1_170 =>
            next_state <= multiplication_with_reduction_special_prime_1_170;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_171;
            end if;
        when multiplication_with_reduction_special_prime_1_171 =>
            next_state <= multiplication_with_reduction_special_prime_1_171;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_172;
            end if;
        when multiplication_with_reduction_special_prime_1_172 =>
            next_state <= multiplication_with_reduction_special_prime_1_172;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_173;
            end if;
        when multiplication_with_reduction_special_prime_1_173 =>
            next_state <= multiplication_with_reduction_special_prime_1_173;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_174;
            end if;
        when multiplication_with_reduction_special_prime_1_174 =>
            next_state <= multiplication_with_reduction_special_prime_1_174;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_175;
            end if;
        when multiplication_with_reduction_special_prime_1_175 =>
            next_state <= multiplication_with_reduction_special_prime_1_175;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_176;
            end if;
        when multiplication_with_reduction_special_prime_1_176 =>
            next_state <= multiplication_with_reduction_special_prime_1_176;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_177;
            end if;
        when multiplication_with_reduction_special_prime_1_177 =>
            next_state <= multiplication_with_reduction_special_prime_1_177;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_178;
            end if;
        when multiplication_with_reduction_special_prime_1_178 =>
            next_state <= multiplication_with_reduction_special_prime_1_178;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_179;
            end if;
        when multiplication_with_reduction_special_prime_1_179 =>
            next_state <= multiplication_with_reduction_special_prime_1_179;
            if(ultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when multiplication_with_reduction_special_prime_1_181 =>
            next_state <= multiplication_with_reduction_special_prime_1_181;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_182;
            end if;
        when multiplication_with_reduction_special_prime_1_182 =>
            next_state <= multiplication_with_reduction_special_prime_1_182;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_183;
            end if;
        when multiplication_with_reduction_special_prime_1_183 =>
            next_state <= multiplication_with_reduction_special_prime_1_183;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_184;
            end if;
        when multiplication_with_reduction_special_prime_1_184 =>
            next_state <= multiplication_with_reduction_special_prime_1_184;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_185;
            end if;
        when multiplication_with_reduction_special_prime_1_185 =>
            next_state <= multiplication_with_reduction_special_prime_1_185;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_186;
            end if;
        when multiplication_with_reduction_special_prime_1_186 =>
            next_state <= multiplication_with_reduction_special_prime_1_186;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_187;
            end if;
        when multiplication_with_reduction_special_prime_1_187 =>
            next_state <= multiplication_with_reduction_special_prime_1_187;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_188;
            end if;
        when multiplication_with_reduction_special_prime_1_188 =>
            next_state <= multiplication_with_reduction_special_prime_1_188;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_189;
            end if;
        when multiplication_with_reduction_special_prime_1_189 =>
            next_state <= multiplication_with_reduction_special_prime_1_189;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_190;
            end if;
        when multiplication_with_reduction_special_prime_1_190 =>
            next_state <= multiplication_with_reduction_special_prime_1_190;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_191;
            end if;
        when multiplication_with_reduction_special_prime_1_191 =>
            next_state <= multiplication_with_reduction_special_prime_1_191;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_192;
            end if;
        when multiplication_with_reduction_special_prime_1_192 =>
            next_state <= multiplication_with_reduction_special_prime_1_192;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_193;
            end if;
        when multiplication_with_reduction_special_prime_1_193 =>
            next_state <= multiplication_with_reduction_special_prime_1_193;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_194;
            end if;
        when multiplication_with_reduction_special_prime_1_194 =>
            next_state <= multiplication_with_reduction_special_prime_1_194;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_195;
            end if;
        when multiplication_with_reduction_special_prime_1_195 =>
            next_state <= multiplication_with_reduction_special_prime_1_195;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_196;
            end if;
        when multiplication_with_reduction_special_prime_1_196 =>
            next_state <= multiplication_with_reduction_special_prime_1_196;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_197;
            end if;
        when multiplication_with_reduction_special_prime_1_197 =>
            next_state <= multiplication_with_reduction_special_prime_1_197;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_198;
            end if;
        when multiplication_with_reduction_special_prime_1_198 =>
            next_state <= multiplication_with_reduction_special_prime_1_198;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_199;
            end if;
        when multiplication_with_reduction_special_prime_1_199 =>
            next_state <= multiplication_with_reduction_special_prime_1_199;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_200;
            end if;
        when multiplication_with_reduction_special_prime_1_200 =>
            next_state <= multiplication_with_reduction_special_prime_1_200;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_201;
            end if;
        when multiplication_with_reduction_special_prime_1_201 =>
            next_state <= multiplication_with_reduction_special_prime_1_201;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_202;
            end if;
        when multiplication_with_reduction_special_prime_1_202 =>
            next_state <= multiplication_with_reduction_special_prime_1_202;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_203;
            end if;
        when multiplication_with_reduction_special_prime_1_203 =>
            next_state <= multiplication_with_reduction_special_prime_1_203;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_204;
            end if;
        when multiplication_with_reduction_special_prime_1_204 =>
            next_state <= multiplication_with_reduction_special_prime_1_204;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_205;
            end if;
        when multiplication_with_reduction_special_prime_1_205 =>
            next_state <= multiplication_with_reduction_special_prime_1_205;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_206;
            end if;
        when multiplication_with_reduction_special_prime_1_206 =>
            next_state <= multiplication_with_reduction_special_prime_1_206;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_207;
            end if;
        when multiplication_with_reduction_special_prime_1_207 =>
            next_state <= multiplication_with_reduction_special_prime_1_207;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_208;
            end if;
        when multiplication_with_reduction_special_prime_1_208 =>
            next_state <= multiplication_with_reduction_special_prime_1_208;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_209;
            end if;
        when multiplication_with_reduction_special_prime_1_209 =>
            next_state <= multiplication_with_reduction_special_prime_1_209;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_210;
            end if;
        when multiplication_with_reduction_special_prime_1_210 =>
            next_state <= multiplication_with_reduction_special_prime_1_210;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_211;
            end if;
        when multiplication_with_reduction_special_prime_1_211 =>
            next_state <= multiplication_with_reduction_special_prime_1_211;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_212;
            end if;
        when multiplication_with_reduction_special_prime_1_212 =>
            next_state <= multiplication_with_reduction_special_prime_1_212;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_213;
            end if;
        when multiplication_with_reduction_special_prime_1_213 =>
            next_state <= multiplication_with_reduction_special_prime_1_213;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_214;
            end if;
        when multiplication_with_reduction_special_prime_1_214 =>
            next_state <= multiplication_with_reduction_special_prime_1_214;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_215;
            end if;
        when multiplication_with_reduction_special_prime_1_215 =>
            next_state <= multiplication_with_reduction_special_prime_1_215;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_216;
            end if;
        when multiplication_with_reduction_special_prime_1_216 =>
            next_state <= multiplication_with_reduction_special_prime_1_216;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_217;
            end if;
        when multiplication_with_reduction_special_prime_1_217 =>
            next_state <= multiplication_with_reduction_special_prime_1_217;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_218;
            end if;
        when multiplication_with_reduction_special_prime_1_218 =>
            next_state <= multiplication_with_reduction_special_prime_1_218;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_219;
            end if;
        when multiplication_with_reduction_special_prime_1_219 =>
            next_state <= multiplication_with_reduction_special_prime_1_219;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_220;
            end if;
        when multiplication_with_reduction_special_prime_1_220 =>
            next_state <= multiplication_with_reduction_special_prime_1_220;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_221;
            end if;
        when multiplication_with_reduction_special_prime_1_221 =>
            next_state <= multiplication_with_reduction_special_prime_1_221;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_222;
            end if;
        when multiplication_with_reduction_special_prime_1_222 =>
            next_state <= multiplication_with_reduction_special_prime_1_222;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_223;
            end if;
        when multiplication_with_reduction_special_prime_1_223 =>
            next_state <= multiplication_with_reduction_special_prime_1_223;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_224;
            end if;
        when multiplication_with_reduction_special_prime_1_224 =>
            next_state <= multiplication_with_reduction_special_prime_1_224;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_225;
            end if;
        when multiplication_with_reduction_special_prime_1_225 =>
            next_state <= multiplication_with_reduction_special_prime_1_225;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_226;
            end if;
        when multiplication_with_reduction_special_prime_1_226 =>
            next_state <= multiplication_with_reduction_special_prime_1_226;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_227;
            end if;
        when multiplication_with_reduction_special_prime_1_227 =>
            next_state <= multiplication_with_reduction_special_prime_1_227;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_228;
            end if;
        when multiplication_with_reduction_special_prime_1_228 =>
            next_state <= multiplication_with_reduction_special_prime_1_228;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_229;
            end if;
        when multiplication_with_reduction_special_prime_1_229 =>
            next_state <= multiplication_with_reduction_special_prime_1_229;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_230;
            end if;
        when multiplication_with_reduction_special_prime_1_230 =>
            next_state <= multiplication_with_reduction_special_prime_1_230;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_231;
            end if;
        when multiplication_with_reduction_special_prime_1_231 =>
            next_state <= multiplication_with_reduction_special_prime_1_231;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_232;
            end if;
        when multiplication_with_reduction_special_prime_1_232 =>
            next_state <= multiplication_with_reduction_special_prime_1_232;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_233;
            end if;
        when multiplication_with_reduction_special_prime_1_233 =>
            next_state <= multiplication_with_reduction_special_prime_1_233;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_234;
            end if;
        when multiplication_with_reduction_special_prime_1_234 =>
            next_state <= multiplication_with_reduction_special_prime_1_234;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_235;
            end if;
        when multiplication_with_reduction_special_prime_1_235 =>
            next_state <= multiplication_with_reduction_special_prime_1_235;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_236;
            end if;
        when multiplication_with_reduction_special_prime_1_236 =>
            next_state <= multiplication_with_reduction_special_prime_1_236;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_237;
            end if;
        when multiplication_with_reduction_special_prime_1_237 =>
            next_state <= multiplication_with_reduction_special_prime_1_237;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_238;
            end if;
        when multiplication_with_reduction_special_prime_1_238 =>
            next_state <= multiplication_with_reduction_special_prime_1_238;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_239;
            end if;
        when multiplication_with_reduction_special_prime_1_239 =>
            next_state <= multiplication_with_reduction_special_prime_1_239;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_240;
            end if;
        when multiplication_with_reduction_special_prime_1_240 =>
            next_state <= multiplication_with_reduction_special_prime_1_240;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_241;
            end if;
        when multiplication_with_reduction_special_prime_1_241 =>
            next_state <= multiplication_with_reduction_special_prime_1_241;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_242;
            end if;
        when multiplication_with_reduction_special_prime_1_242 =>
            next_state <= multiplication_with_reduction_special_prime_1_242;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_243;
            end if;
        when multiplication_with_reduction_special_prime_1_243 =>
            next_state <= multiplication_with_reduction_special_prime_1_243;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_244;
            end if;
        when multiplication_with_reduction_special_prime_1_244 =>
            next_state <= multiplication_with_reduction_special_prime_1_244;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_245;
            end if;
        when multiplication_with_reduction_special_prime_1_245 =>
            next_state <= multiplication_with_reduction_special_prime_1_245;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_246;
            end if;
        when multiplication_with_reduction_special_prime_1_246 =>
            next_state <= multiplication_with_reduction_special_prime_1_246;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_247;
            end if;
        when multiplication_with_reduction_special_prime_1_247 =>
            next_state <= multiplication_with_reduction_special_prime_1_247;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_248;
            end if;
        when multiplication_with_reduction_special_prime_1_248 =>
            next_state <= multiplication_with_reduction_special_prime_1_248;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_249;
            end if;
        when multiplication_with_reduction_special_prime_1_249 =>
            next_state <= multiplication_with_reduction_special_prime_1_249;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_250;
            end if;
        when multiplication_with_reduction_special_prime_1_250 =>
            next_state <= multiplication_with_reduction_special_prime_1_250;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_251;
            end if;
        when multiplication_with_reduction_special_prime_1_251 =>
            next_state <= multiplication_with_reduction_special_prime_1_251;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_252;
            end if;
        when multiplication_with_reduction_special_prime_1_252 =>
            next_state <= multiplication_with_reduction_special_prime_1_252;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1_253;
            end if;
        when multiplication_with_reduction_special_prime_1_253 =>
            next_state <= multiplication_with_reduction_special_prime_1_253;
            if(ultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when multiplication_with_reduction_special_prime_2_0 => 
            next_state <= multiplication_with_reduction_special_prime_2_0;
            if(ultimate_operation = '1') then
                if(operands_size = "001") then
                    next_state <= multiplication_with_reduction_special_prime_2_1;
                else
                    next_state <= multiplication_with_reduction_special_prime_2_5;
                end if;
            end if;
        when multiplication_with_reduction_special_prime_2_1 => 
            next_state <= multiplication_with_reduction_special_prime_2_1;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_2;
            end if;
        when multiplication_with_reduction_special_prime_2_2 => 
            next_state <= multiplication_with_reduction_special_prime_2_2;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_3;
            end if;
        when multiplication_with_reduction_special_prime_2_3 => 
            next_state <= multiplication_with_reduction_special_prime_2_3;
            if(ultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when multiplication_with_reduction_special_prime_2_5 => 
            next_state <= multiplication_with_reduction_special_prime_2_5;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_6;
            end if;
        when multiplication_with_reduction_special_prime_2_6 => 
            next_state <= multiplication_with_reduction_special_prime_2_6;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_7;
            end if;
        when multiplication_with_reduction_special_prime_2_7 => 
            next_state <= multiplication_with_reduction_special_prime_2_7;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_8;
            end if;
        when multiplication_with_reduction_special_prime_2_8 => 
            next_state <= multiplication_with_reduction_special_prime_2_8;
            if(ultimate_operation = '1') then
                if(operands_size = "010") then
                    next_state <= multiplication_with_reduction_special_prime_2_9;
                else
                    next_state <= multiplication_with_reduction_special_prime_2_17;
                end if;
            end if;
        when multiplication_with_reduction_special_prime_2_9 => 
            next_state <= multiplication_with_reduction_special_prime_2_9;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_10;
            end if;
        when multiplication_with_reduction_special_prime_2_10 => 
            next_state <= multiplication_with_reduction_special_prime_2_10;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_11;
            end if;
        when multiplication_with_reduction_special_prime_2_11 => 
            next_state <= multiplication_with_reduction_special_prime_2_11;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_12;
            end if;
        when multiplication_with_reduction_special_prime_2_12 => 
            next_state <= multiplication_with_reduction_special_prime_2_12;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_13;
            end if;
        when multiplication_with_reduction_special_prime_2_13 => 
            next_state <= multiplication_with_reduction_special_prime_2_13;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_14;
            end if;
        when multiplication_with_reduction_special_prime_2_14 => 
            next_state <= multiplication_with_reduction_special_prime_2_14;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_15;
            end if;
        when multiplication_with_reduction_special_prime_2_15 => 
            next_state <= multiplication_with_reduction_special_prime_2_15;
            if(ultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when multiplication_with_reduction_special_prime_2_17 => 
            next_state <= multiplication_with_reduction_special_prime_2_17;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_18;
            end if;
        when multiplication_with_reduction_special_prime_2_18 => 
            next_state <= multiplication_with_reduction_special_prime_2_18;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_19;
            end if;
        when multiplication_with_reduction_special_prime_2_19 => 
            next_state <= multiplication_with_reduction_special_prime_2_19;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_20;
            end if;
        when multiplication_with_reduction_special_prime_2_20 => 
            next_state <= multiplication_with_reduction_special_prime_2_20;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_21;
            end if;
        when multiplication_with_reduction_special_prime_2_21 => 
            next_state <= multiplication_with_reduction_special_prime_2_21;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_22;
            end if;
        when multiplication_with_reduction_special_prime_2_22 => 
            next_state <= multiplication_with_reduction_special_prime_2_22;
            if(ultimate_operation = '1') then
                if(operands_size = "011") then
                    next_state <= multiplication_with_reduction_special_prime_2_23;
                else
                    next_state <= multiplication_with_reduction_special_prime_2_37;
                end if;
            end if;
        when multiplication_with_reduction_special_prime_2_23 => 
            next_state <= multiplication_with_reduction_special_prime_2_23;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_24;
            end if;
        when multiplication_with_reduction_special_prime_2_24 => 
            next_state <= multiplication_with_reduction_special_prime_2_24;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_25;
            end if;
        when multiplication_with_reduction_special_prime_2_25 => 
            next_state <= multiplication_with_reduction_special_prime_2_25;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_26;
            end if;
        when multiplication_with_reduction_special_prime_2_26 => 
            next_state <= multiplication_with_reduction_special_prime_2_26;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_27;
            end if;
        when multiplication_with_reduction_special_prime_2_27 => 
            next_state <= multiplication_with_reduction_special_prime_2_27;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_28;
            end if;
        when multiplication_with_reduction_special_prime_2_28 => 
            next_state <= multiplication_with_reduction_special_prime_2_28;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_29;
            end if;
        when multiplication_with_reduction_special_prime_2_29 => 
            next_state <= multiplication_with_reduction_special_prime_2_29;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_30;
            end if;
        when multiplication_with_reduction_special_prime_2_30 => 
            next_state <= multiplication_with_reduction_special_prime_2_30;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_31;
            end if;
        when multiplication_with_reduction_special_prime_2_31 => 
            next_state <= multiplication_with_reduction_special_prime_2_31;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_32;
            end if;
        when multiplication_with_reduction_special_prime_2_32 => 
            next_state <= multiplication_with_reduction_special_prime_2_32;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_33;
            end if;
        when multiplication_with_reduction_special_prime_2_33 => 
            next_state <= multiplication_with_reduction_special_prime_2_33;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_34;
            end if;
        when multiplication_with_reduction_special_prime_2_34 => 
            next_state <= multiplication_with_reduction_special_prime_2_34;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_35;
            end if;
        when multiplication_with_reduction_special_prime_2_35 => 
            next_state <= multiplication_with_reduction_special_prime_2_35;
            if(ultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when multiplication_with_reduction_special_prime_2_37 => 
            next_state <= multiplication_with_reduction_special_prime_2_37;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_38;
            end if;
        when multiplication_with_reduction_special_prime_2_38 => 
            next_state <= multiplication_with_reduction_special_prime_2_38;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_39;
            end if;
        when multiplication_with_reduction_special_prime_2_39 => 
            next_state <= multiplication_with_reduction_special_prime_2_39;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_40;
            end if;
        when multiplication_with_reduction_special_prime_2_40 => 
            next_state <= multiplication_with_reduction_special_prime_2_40;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_41;
            end if;
        when multiplication_with_reduction_special_prime_2_41 => 
            next_state <= multiplication_with_reduction_special_prime_2_41;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_42;
            end if;
        when multiplication_with_reduction_special_prime_2_42 => 
            next_state <= multiplication_with_reduction_special_prime_2_42;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_43;
            end if;
        when multiplication_with_reduction_special_prime_2_43 => 
            next_state <= multiplication_with_reduction_special_prime_2_43;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_44;
            end if;
        when multiplication_with_reduction_special_prime_2_44 => 
            next_state <= multiplication_with_reduction_special_prime_2_44;
            if(ultimate_operation = '1') then
                if(operands_size = "100") then
                    next_state <= multiplication_with_reduction_special_prime_2_45;
                else
                    next_state <= multiplication_with_reduction_special_prime_2_67;
                end if;
            end if;
        when multiplication_with_reduction_special_prime_2_45 => 
            next_state <= multiplication_with_reduction_special_prime_2_45;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_46;
            end if;
        when multiplication_with_reduction_special_prime_2_46 => 
            next_state <= multiplication_with_reduction_special_prime_2_46;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_47;
            end if;
        when multiplication_with_reduction_special_prime_2_47 => 
            next_state <= multiplication_with_reduction_special_prime_2_47;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_48;
            end if;
        when multiplication_with_reduction_special_prime_2_48 => 
            next_state <= multiplication_with_reduction_special_prime_2_48;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_49;
            end if;
        when multiplication_with_reduction_special_prime_2_49 => 
            next_state <= multiplication_with_reduction_special_prime_2_49;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_50;
            end if;
        when multiplication_with_reduction_special_prime_2_50 => 
            next_state <= multiplication_with_reduction_special_prime_2_50;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_51;
            end if;
        when multiplication_with_reduction_special_prime_2_51 => 
            next_state <= multiplication_with_reduction_special_prime_2_51;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_52;
            end if;
        when multiplication_with_reduction_special_prime_2_52 => 
            next_state <= multiplication_with_reduction_special_prime_2_52;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_53;
            end if;
        when multiplication_with_reduction_special_prime_2_53 => 
            next_state <= multiplication_with_reduction_special_prime_2_53;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_54;
            end if;
        when multiplication_with_reduction_special_prime_2_54 => 
            next_state <= multiplication_with_reduction_special_prime_2_54;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_55;
            end if;
        when multiplication_with_reduction_special_prime_2_55 => 
            next_state <= multiplication_with_reduction_special_prime_2_55;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_56;
            end if;
        when multiplication_with_reduction_special_prime_2_56 => 
            next_state <= multiplication_with_reduction_special_prime_2_56;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_57;
            end if;
        when multiplication_with_reduction_special_prime_2_57 => 
            next_state <= multiplication_with_reduction_special_prime_2_57;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_58;
            end if;
        when multiplication_with_reduction_special_prime_2_58 => 
            next_state <= multiplication_with_reduction_special_prime_2_58;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_59;
            end if;
        when multiplication_with_reduction_special_prime_2_59 => 
            next_state <= multiplication_with_reduction_special_prime_2_59;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_60;
            end if;
        when multiplication_with_reduction_special_prime_2_60 => 
            next_state <= multiplication_with_reduction_special_prime_2_60;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_61;
            end if;
        when multiplication_with_reduction_special_prime_2_61 => 
            next_state <= multiplication_with_reduction_special_prime_2_61;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_62;
            end if;
        when multiplication_with_reduction_special_prime_2_62 => 
            next_state <= multiplication_with_reduction_special_prime_2_62;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_63;
            end if;
        when multiplication_with_reduction_special_prime_2_63 => 
            next_state <= multiplication_with_reduction_special_prime_2_63;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_64;
            end if;
        when multiplication_with_reduction_special_prime_2_64 => 
            next_state <= multiplication_with_reduction_special_prime_2_64;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_65;
            end if;
        when multiplication_with_reduction_special_prime_2_65 => 
            next_state <= multiplication_with_reduction_special_prime_2_65;
            if(ultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when multiplication_with_reduction_special_prime_2_67 => 
            next_state <= multiplication_with_reduction_special_prime_2_67;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_68;
            end if;
        when multiplication_with_reduction_special_prime_2_68 => 
            next_state <= multiplication_with_reduction_special_prime_2_68;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_69;
            end if;
        when multiplication_with_reduction_special_prime_2_69 => 
            next_state <= multiplication_with_reduction_special_prime_2_69;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_70;
            end if;
        when multiplication_with_reduction_special_prime_2_70 => 
            next_state <= multiplication_with_reduction_special_prime_2_70;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_71;
            end if;
        when multiplication_with_reduction_special_prime_2_71 => 
            next_state <= multiplication_with_reduction_special_prime_2_71;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_72;
            end if;
        when multiplication_with_reduction_special_prime_2_72 => 
            next_state <= multiplication_with_reduction_special_prime_2_72;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_73;
            end if;
        when multiplication_with_reduction_special_prime_2_73 => 
            next_state <= multiplication_with_reduction_special_prime_2_73;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_74;
            end if;
        when multiplication_with_reduction_special_prime_2_74 => 
            next_state <= multiplication_with_reduction_special_prime_2_74;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_75;
            end if;
        when multiplication_with_reduction_special_prime_2_75 => 
            next_state <= multiplication_with_reduction_special_prime_2_75;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_76;
            end if;
        when multiplication_with_reduction_special_prime_2_76 => 
            next_state <= multiplication_with_reduction_special_prime_2_76;
            if(ultimate_operation = '1') then
                if(operands_size = "101") then
                    next_state <= multiplication_with_reduction_special_prime_2_77;
                else
                    next_state <= multiplication_with_reduction_special_prime_2_109;
                end if;
            end if;
        when multiplication_with_reduction_special_prime_2_77 => 
            next_state <= multiplication_with_reduction_special_prime_2_77;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_78;
            end if;
        when multiplication_with_reduction_special_prime_2_78 => 
            next_state <= multiplication_with_reduction_special_prime_2_78;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_79;
            end if;
        when multiplication_with_reduction_special_prime_2_79 => 
            next_state <= multiplication_with_reduction_special_prime_2_79;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_80;
            end if;
        when multiplication_with_reduction_special_prime_2_80 => 
            next_state <= multiplication_with_reduction_special_prime_2_80;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_81;
            end if;
        when multiplication_with_reduction_special_prime_2_81 => 
            next_state <= multiplication_with_reduction_special_prime_2_81;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_82;
            end if;
        when multiplication_with_reduction_special_prime_2_82 => 
            next_state <= multiplication_with_reduction_special_prime_2_82;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_83;
            end if;
        when multiplication_with_reduction_special_prime_2_83 => 
            next_state <= multiplication_with_reduction_special_prime_2_83;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_84;
            end if;
        when multiplication_with_reduction_special_prime_2_84 => 
            next_state <= multiplication_with_reduction_special_prime_2_84;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_85;
            end if;
        when multiplication_with_reduction_special_prime_2_85 => 
            next_state <= multiplication_with_reduction_special_prime_2_85;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_86;
            end if;
        when multiplication_with_reduction_special_prime_2_86 => 
            next_state <= multiplication_with_reduction_special_prime_2_86;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_87;
            end if;
        when multiplication_with_reduction_special_prime_2_87 => 
            next_state <= multiplication_with_reduction_special_prime_2_87;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_88;
            end if;
        when multiplication_with_reduction_special_prime_2_88 => 
            next_state <= multiplication_with_reduction_special_prime_2_88;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_89;
            end if;
        when multiplication_with_reduction_special_prime_2_89 => 
            next_state <= multiplication_with_reduction_special_prime_2_89;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_90;
            end if;
        when multiplication_with_reduction_special_prime_2_90 => 
            next_state <= multiplication_with_reduction_special_prime_2_90;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_91;
            end if;
        when multiplication_with_reduction_special_prime_2_91 => 
            next_state <= multiplication_with_reduction_special_prime_2_91;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_92;
            end if;
        when multiplication_with_reduction_special_prime_2_92 => 
            next_state <= multiplication_with_reduction_special_prime_2_92;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_93;
            end if;
        when multiplication_with_reduction_special_prime_2_93 => 
            next_state <= multiplication_with_reduction_special_prime_2_93;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_94;
            end if;
        when multiplication_with_reduction_special_prime_2_94 => 
            next_state <= multiplication_with_reduction_special_prime_2_94;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_95;
            end if;
        when multiplication_with_reduction_special_prime_2_95 => 
            next_state <= multiplication_with_reduction_special_prime_2_95;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_96;
            end if;
        when multiplication_with_reduction_special_prime_2_96 => 
            next_state <= multiplication_with_reduction_special_prime_2_96;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_97;
            end if;
        when multiplication_with_reduction_special_prime_2_97 => 
            next_state <= multiplication_with_reduction_special_prime_2_97;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_98;
            end if;
        when multiplication_with_reduction_special_prime_2_98 => 
            next_state <= multiplication_with_reduction_special_prime_2_98;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_99;
            end if;
        when multiplication_with_reduction_special_prime_2_99 => 
            next_state <= multiplication_with_reduction_special_prime_2_99;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_100;
            end if;
        when multiplication_with_reduction_special_prime_2_100 => 
            next_state <= multiplication_with_reduction_special_prime_2_100;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_101;
            end if;
        when multiplication_with_reduction_special_prime_2_101 => 
            next_state <= multiplication_with_reduction_special_prime_2_101;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_102;
            end if;
        when multiplication_with_reduction_special_prime_2_102 => 
            next_state <= multiplication_with_reduction_special_prime_2_102;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_103;
            end if;
        when multiplication_with_reduction_special_prime_2_103 => 
            next_state <= multiplication_with_reduction_special_prime_2_103;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_104;
            end if;
        when multiplication_with_reduction_special_prime_2_104 => 
            next_state <= multiplication_with_reduction_special_prime_2_104;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_105;
            end if;
        when multiplication_with_reduction_special_prime_2_105 => 
            next_state <= multiplication_with_reduction_special_prime_2_105;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_106;
            end if;
        when multiplication_with_reduction_special_prime_2_106 => 
            next_state <= multiplication_with_reduction_special_prime_2_106;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_107;
            end if;
        when multiplication_with_reduction_special_prime_2_107 => 
            next_state <= multiplication_with_reduction_special_prime_2_107;
            if(ultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when multiplication_with_reduction_special_prime_2_109 => 
            next_state <= multiplication_with_reduction_special_prime_2_109;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_110;
            end if;
        when multiplication_with_reduction_special_prime_2_110 => 
            next_state <= multiplication_with_reduction_special_prime_2_110;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_111;
            end if;
        when multiplication_with_reduction_special_prime_2_111 => 
            next_state <= multiplication_with_reduction_special_prime_2_111;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_112;
            end if;
        when multiplication_with_reduction_special_prime_2_112 => 
            next_state <= multiplication_with_reduction_special_prime_2_112;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_113;
            end if;
        when multiplication_with_reduction_special_prime_2_113 => 
            next_state <= multiplication_with_reduction_special_prime_2_113;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_114;
            end if;
        when multiplication_with_reduction_special_prime_2_114 => 
            next_state <= multiplication_with_reduction_special_prime_2_114;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_115;
            end if;
        when multiplication_with_reduction_special_prime_2_115 => 
            next_state <= multiplication_with_reduction_special_prime_2_115;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_116;
            end if;
        when multiplication_with_reduction_special_prime_2_116 => 
            next_state <= multiplication_with_reduction_special_prime_2_116;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_117;
            end if;
        when multiplication_with_reduction_special_prime_2_117 => 
            next_state <= multiplication_with_reduction_special_prime_2_117;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_118;
            end if;
        when multiplication_with_reduction_special_prime_2_118 => 
            next_state <= multiplication_with_reduction_special_prime_2_118;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_119;
            end if;
        when multiplication_with_reduction_special_prime_2_119 => 
            next_state <= multiplication_with_reduction_special_prime_2_119;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_120;
            end if;
        when multiplication_with_reduction_special_prime_2_120 => 
            next_state <= multiplication_with_reduction_special_prime_2_120;
            if(ultimate_operation = '1') then
                if(operands_size = "110") then
                    next_state <= multiplication_with_reduction_special_prime_2_121;
                else
                    next_state <= multiplication_with_reduction_special_prime_2_165;
                end if;
            end if;
        when multiplication_with_reduction_special_prime_2_121 => 
            next_state <= multiplication_with_reduction_special_prime_2_121;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_122;
            end if;
        when multiplication_with_reduction_special_prime_2_122 => 
            next_state <= multiplication_with_reduction_special_prime_2_122;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_123;
            end if;
        when multiplication_with_reduction_special_prime_2_123 => 
            next_state <= multiplication_with_reduction_special_prime_2_123;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_124;
            end if;
        when multiplication_with_reduction_special_prime_2_124 => 
            next_state <= multiplication_with_reduction_special_prime_2_124;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_125;
            end if;
        when multiplication_with_reduction_special_prime_2_125 => 
            next_state <= multiplication_with_reduction_special_prime_2_125;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_126;
            end if;
        when multiplication_with_reduction_special_prime_2_126 => 
            next_state <= multiplication_with_reduction_special_prime_2_126;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_127;
            end if;
        when multiplication_with_reduction_special_prime_2_127 => 
            next_state <= multiplication_with_reduction_special_prime_2_127;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_128;
            end if;
        when multiplication_with_reduction_special_prime_2_128 => 
            next_state <= multiplication_with_reduction_special_prime_2_128;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_129;
            end if;
        when multiplication_with_reduction_special_prime_2_129 => 
            next_state <= multiplication_with_reduction_special_prime_2_129;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_130;
            end if;
        when multiplication_with_reduction_special_prime_2_130 => 
            next_state <= multiplication_with_reduction_special_prime_2_130;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_131;
            end if;
        when multiplication_with_reduction_special_prime_2_131 => 
            next_state <= multiplication_with_reduction_special_prime_2_131;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_132;
            end if;
        when multiplication_with_reduction_special_prime_2_132 => 
            next_state <= multiplication_with_reduction_special_prime_2_132;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_133;
            end if;
        when multiplication_with_reduction_special_prime_2_133 => 
            next_state <= multiplication_with_reduction_special_prime_2_133;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_134;
            end if;
        when multiplication_with_reduction_special_prime_2_134 => 
            next_state <= multiplication_with_reduction_special_prime_2_134;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_135;
            end if;
        when multiplication_with_reduction_special_prime_2_135 => 
            next_state <= multiplication_with_reduction_special_prime_2_135;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_136;
            end if;
        when multiplication_with_reduction_special_prime_2_136 => 
            next_state <= multiplication_with_reduction_special_prime_2_136;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_137;
            end if;
        when multiplication_with_reduction_special_prime_2_137 => 
            next_state <= multiplication_with_reduction_special_prime_2_137;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_138;
            end if;
        when multiplication_with_reduction_special_prime_2_138 => 
            next_state <= multiplication_with_reduction_special_prime_2_138;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_139;
            end if;
        when multiplication_with_reduction_special_prime_2_139 => 
            next_state <= multiplication_with_reduction_special_prime_2_139;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_140;
            end if;
        when multiplication_with_reduction_special_prime_2_140 => 
            next_state <= multiplication_with_reduction_special_prime_2_140;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_141;
            end if;
        when multiplication_with_reduction_special_prime_2_141 => 
            next_state <= multiplication_with_reduction_special_prime_2_141;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_142;
            end if;
        when multiplication_with_reduction_special_prime_2_142 => 
            next_state <= multiplication_with_reduction_special_prime_2_142;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_143;
            end if;
        when multiplication_with_reduction_special_prime_2_143 => 
            next_state <= multiplication_with_reduction_special_prime_2_143;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_144;
            end if;
        when multiplication_with_reduction_special_prime_2_144 => 
            next_state <= multiplication_with_reduction_special_prime_2_144;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_145;
            end if;
        when multiplication_with_reduction_special_prime_2_145 => 
            next_state <= multiplication_with_reduction_special_prime_2_145;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_146;
            end if;
        when multiplication_with_reduction_special_prime_2_146 => 
            next_state <= multiplication_with_reduction_special_prime_2_146;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_147;
            end if;
        when multiplication_with_reduction_special_prime_2_147 => 
            next_state <= multiplication_with_reduction_special_prime_2_147;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_148;
            end if;
        when multiplication_with_reduction_special_prime_2_148 => 
            next_state <= multiplication_with_reduction_special_prime_2_148;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_149;
            end if;
        when multiplication_with_reduction_special_prime_2_149 => 
            next_state <= multiplication_with_reduction_special_prime_2_149;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_150;
            end if;
        when multiplication_with_reduction_special_prime_2_150 => 
            next_state <= multiplication_with_reduction_special_prime_2_150;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_151;
            end if;
        when multiplication_with_reduction_special_prime_2_151 => 
            next_state <= multiplication_with_reduction_special_prime_2_151;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_152;
            end if;
        when multiplication_with_reduction_special_prime_2_152 => 
            next_state <= multiplication_with_reduction_special_prime_2_152;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_153;
            end if;
        when multiplication_with_reduction_special_prime_2_153 => 
            next_state <= multiplication_with_reduction_special_prime_2_153;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_154;
            end if;
        when multiplication_with_reduction_special_prime_2_154 => 
            next_state <= multiplication_with_reduction_special_prime_2_154;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_155;
            end if;
        when multiplication_with_reduction_special_prime_2_155 => 
            next_state <= multiplication_with_reduction_special_prime_2_155;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_156;
            end if;
        when multiplication_with_reduction_special_prime_2_156 => 
            next_state <= multiplication_with_reduction_special_prime_2_156;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_157;
            end if;
        when multiplication_with_reduction_special_prime_2_157 => 
            next_state <= multiplication_with_reduction_special_prime_2_157;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_158;
            end if;
        when multiplication_with_reduction_special_prime_2_158 => 
            next_state <= multiplication_with_reduction_special_prime_2_158;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_159;
            end if;
        when multiplication_with_reduction_special_prime_2_159 => 
            next_state <= multiplication_with_reduction_special_prime_2_159;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_160;
            end if;
        when multiplication_with_reduction_special_prime_2_160 => 
            next_state <= multiplication_with_reduction_special_prime_2_160;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_161;
            end if;
        when multiplication_with_reduction_special_prime_2_161 => 
            next_state <= multiplication_with_reduction_special_prime_2_161;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_162;
            end if;
        when multiplication_with_reduction_special_prime_2_162 => 
            next_state <= multiplication_with_reduction_special_prime_2_162;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_163;
            end if;
        when multiplication_with_reduction_special_prime_2_163 => 
            next_state <= multiplication_with_reduction_special_prime_2_163;
            if(ultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when multiplication_with_reduction_special_prime_2_165 => 
            next_state <= multiplication_with_reduction_special_prime_2_165;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_166;
            end if;
        when multiplication_with_reduction_special_prime_2_166 => 
            next_state <= multiplication_with_reduction_special_prime_2_166;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_167;
            end if;
        when multiplication_with_reduction_special_prime_2_167 => 
            next_state <= multiplication_with_reduction_special_prime_2_167;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_168;
            end if;
        when multiplication_with_reduction_special_prime_2_168 => 
            next_state <= multiplication_with_reduction_special_prime_2_168;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_169;
            end if;
        when multiplication_with_reduction_special_prime_2_169 => 
            next_state <= multiplication_with_reduction_special_prime_2_169;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_170;
            end if;
        when multiplication_with_reduction_special_prime_2_170 => 
            next_state <= multiplication_with_reduction_special_prime_2_170;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_171;
            end if;
        when multiplication_with_reduction_special_prime_2_171 => 
            next_state <= multiplication_with_reduction_special_prime_2_171;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_172;
            end if;
        when multiplication_with_reduction_special_prime_2_172 => 
            next_state <= multiplication_with_reduction_special_prime_2_172;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_173;
            end if;
        when multiplication_with_reduction_special_prime_2_173 => 
            next_state <= multiplication_with_reduction_special_prime_2_173;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_174;
            end if;
        when multiplication_with_reduction_special_prime_2_174 => 
            next_state <= multiplication_with_reduction_special_prime_2_174;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_175;
            end if;
        when multiplication_with_reduction_special_prime_2_175 => 
            next_state <= multiplication_with_reduction_special_prime_2_175;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_176;
            end if;
        when multiplication_with_reduction_special_prime_2_176 => 
            next_state <= multiplication_with_reduction_special_prime_2_176;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_177;
            end if;
        when multiplication_with_reduction_special_prime_2_177 => 
            next_state <= multiplication_with_reduction_special_prime_2_177;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_178;
            end if;
        when multiplication_with_reduction_special_prime_2_178 => 
            next_state <= multiplication_with_reduction_special_prime_2_178;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_179;
            end if;
        when multiplication_with_reduction_special_prime_2_179 => 
            next_state <= multiplication_with_reduction_special_prime_2_179;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_180;
            end if;
        when multiplication_with_reduction_special_prime_2_180 => 
            next_state <= multiplication_with_reduction_special_prime_2_180;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_181;
            end if;
        when multiplication_with_reduction_special_prime_2_181 => 
            next_state <= multiplication_with_reduction_special_prime_2_181;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_182;
            end if;
        when multiplication_with_reduction_special_prime_2_182 => 
            next_state <= multiplication_with_reduction_special_prime_2_182;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_183;
            end if;
        when multiplication_with_reduction_special_prime_2_183 => 
            next_state <= multiplication_with_reduction_special_prime_2_183;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_184;
            end if;
        when multiplication_with_reduction_special_prime_2_184 => 
            next_state <= multiplication_with_reduction_special_prime_2_184;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_185;
            end if;
        when multiplication_with_reduction_special_prime_2_185 => 
            next_state <= multiplication_with_reduction_special_prime_2_185;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_186;
            end if;
        when multiplication_with_reduction_special_prime_2_186 => 
            next_state <= multiplication_with_reduction_special_prime_2_186;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_187;
            end if;
        when multiplication_with_reduction_special_prime_2_187 => 
            next_state <= multiplication_with_reduction_special_prime_2_187;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_188;
            end if;
        when multiplication_with_reduction_special_prime_2_188 => 
            next_state <= multiplication_with_reduction_special_prime_2_188;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_189;
            end if;
        when multiplication_with_reduction_special_prime_2_189 => 
            next_state <= multiplication_with_reduction_special_prime_2_189;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_190;
            end if;
        when multiplication_with_reduction_special_prime_2_190 => 
            next_state <= multiplication_with_reduction_special_prime_2_190;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_191;
            end if;
        when multiplication_with_reduction_special_prime_2_191 => 
            next_state <= multiplication_with_reduction_special_prime_2_191;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_192;
            end if;
        when multiplication_with_reduction_special_prime_2_192 => 
            next_state <= multiplication_with_reduction_special_prime_2_192;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_193;
            end if;
        when multiplication_with_reduction_special_prime_2_193 => 
            next_state <= multiplication_with_reduction_special_prime_2_193;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_194;
            end if;
        when multiplication_with_reduction_special_prime_2_194 => 
            next_state <= multiplication_with_reduction_special_prime_2_194;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_195;
            end if;
        when multiplication_with_reduction_special_prime_2_195 => 
            next_state <= multiplication_with_reduction_special_prime_2_195;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_196;
            end if;
        when multiplication_with_reduction_special_prime_2_196 => 
            next_state <= multiplication_with_reduction_special_prime_2_196;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_197;
            end if;
        when multiplication_with_reduction_special_prime_2_197 => 
            next_state <= multiplication_with_reduction_special_prime_2_197;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_198;
            end if;
        when multiplication_with_reduction_special_prime_2_198 => 
            next_state <= multiplication_with_reduction_special_prime_2_198;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_199;
            end if;
        when multiplication_with_reduction_special_prime_2_199 => 
            next_state <= multiplication_with_reduction_special_prime_2_199;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_200;
            end if;
        when multiplication_with_reduction_special_prime_2_200 => 
            next_state <= multiplication_with_reduction_special_prime_2_200;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_201;
            end if;
        when multiplication_with_reduction_special_prime_2_201 => 
            next_state <= multiplication_with_reduction_special_prime_2_201;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_202;
            end if;
        when multiplication_with_reduction_special_prime_2_202 => 
            next_state <= multiplication_with_reduction_special_prime_2_202;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_203;
            end if;
        when multiplication_with_reduction_special_prime_2_203 => 
            next_state <= multiplication_with_reduction_special_prime_2_203;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_204;
            end if;
        when multiplication_with_reduction_special_prime_2_204 => 
            next_state <= multiplication_with_reduction_special_prime_2_204;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_205;
            end if;
        when multiplication_with_reduction_special_prime_2_205 => 
            next_state <= multiplication_with_reduction_special_prime_2_205;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_206;
            end if;
        when multiplication_with_reduction_special_prime_2_206 => 
            next_state <= multiplication_with_reduction_special_prime_2_206;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_207;
            end if;
        when multiplication_with_reduction_special_prime_2_207 => 
            next_state <= multiplication_with_reduction_special_prime_2_207;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_208;
            end if;
        when multiplication_with_reduction_special_prime_2_208 => 
            next_state <= multiplication_with_reduction_special_prime_2_208;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_209;
            end if;
        when multiplication_with_reduction_special_prime_2_209 => 
            next_state <= multiplication_with_reduction_special_prime_2_209;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_210;
            end if;
        when multiplication_with_reduction_special_prime_2_210 => 
            next_state <= multiplication_with_reduction_special_prime_2_210;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_211;
            end if;
        when multiplication_with_reduction_special_prime_2_211 => 
            next_state <= multiplication_with_reduction_special_prime_2_211;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_212;
            end if;
        when multiplication_with_reduction_special_prime_2_212 => 
            next_state <= multiplication_with_reduction_special_prime_2_212;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_213;
            end if;
        when multiplication_with_reduction_special_prime_2_213 => 
            next_state <= multiplication_with_reduction_special_prime_2_213;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_214;
            end if;
        when multiplication_with_reduction_special_prime_2_214 => 
            next_state <= multiplication_with_reduction_special_prime_2_214;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_215;
            end if;
        when multiplication_with_reduction_special_prime_2_215 => 
            next_state <= multiplication_with_reduction_special_prime_2_215;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_216;
            end if;
        when multiplication_with_reduction_special_prime_2_216 => 
            next_state <= multiplication_with_reduction_special_prime_2_216;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_217;
            end if;
        when multiplication_with_reduction_special_prime_2_217 => 
            next_state <= multiplication_with_reduction_special_prime_2_217;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_218;
            end if;
        when multiplication_with_reduction_special_prime_2_218 => 
            next_state <= multiplication_with_reduction_special_prime_2_218;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_219;
            end if;
        when multiplication_with_reduction_special_prime_2_219 => 
            next_state <= multiplication_with_reduction_special_prime_2_219;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_220;
            end if;
        when multiplication_with_reduction_special_prime_2_220 => 
            next_state <= multiplication_with_reduction_special_prime_2_220;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_221;
            end if;
        when multiplication_with_reduction_special_prime_2_221 => 
            next_state <= multiplication_with_reduction_special_prime_2_221;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_222;
            end if;
        when multiplication_with_reduction_special_prime_2_222 => 
            next_state <= multiplication_with_reduction_special_prime_2_222;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_223;
            end if;
        when multiplication_with_reduction_special_prime_2_223 => 
            next_state <= multiplication_with_reduction_special_prime_2_223;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_224;
            end if;
        when multiplication_with_reduction_special_prime_2_224 => 
            next_state <= multiplication_with_reduction_special_prime_2_224;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_225;
            end if;
        when multiplication_with_reduction_special_prime_2_225 => 
            next_state <= multiplication_with_reduction_special_prime_2_225;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_226;
            end if;
        when multiplication_with_reduction_special_prime_2_226 => 
            next_state <= multiplication_with_reduction_special_prime_2_226;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_227;
            end if;
        when multiplication_with_reduction_special_prime_2_227 => 
            next_state <= multiplication_with_reduction_special_prime_2_227;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_228;
            end if;
        when multiplication_with_reduction_special_prime_2_228 => 
            next_state <= multiplication_with_reduction_special_prime_2_228;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_229;
            end if;
        when multiplication_with_reduction_special_prime_2_229 => 
            next_state <= multiplication_with_reduction_special_prime_2_229;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_230;
            end if;
        when multiplication_with_reduction_special_prime_2_230 => 
            next_state <= multiplication_with_reduction_special_prime_2_230;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_231;
            end if;
        when multiplication_with_reduction_special_prime_2_231 => 
            next_state <= multiplication_with_reduction_special_prime_2_231;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_232;
            end if;
        when multiplication_with_reduction_special_prime_2_232 => 
            next_state <= multiplication_with_reduction_special_prime_2_232;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_233;
            end if;
        when multiplication_with_reduction_special_prime_2_233 => 
            next_state <= multiplication_with_reduction_special_prime_2_233;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_234;
            end if;
        when multiplication_with_reduction_special_prime_2_234 => 
            next_state <= multiplication_with_reduction_special_prime_2_234;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_2_235;
            end if;
        when multiplication_with_reduction_special_prime_2_235 => 
            next_state <= multiplication_with_reduction_special_prime_2_235;
            if(ultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when multiplication_with_reduction_special_prime_3_0 =>
            next_state <= multiplication_with_reduction_special_prime_3_0;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_1;
            end if;
        when multiplication_with_reduction_special_prime_3_1 =>
            next_state <= multiplication_with_reduction_special_prime_3_1;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_2;
            end if;
        when multiplication_with_reduction_special_prime_3_2 =>
            next_state <= multiplication_with_reduction_special_prime_3_2;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_3;
            end if;
        when multiplication_with_reduction_special_prime_3_3 =>
            next_state <= multiplication_with_reduction_special_prime_3_3;
            if(ultimate_operation = '1') then
                if(operands_size = "010") then
                    next_state <= multiplication_with_reduction_special_prime_3_4;
                else
                    next_state <= multiplication_with_reduction_special_prime_3_10;
                end if;
            end if;
        when multiplication_with_reduction_special_prime_3_4 =>
            next_state <= multiplication_with_reduction_special_prime_3_4;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_5;
            end if;
        when multiplication_with_reduction_special_prime_3_5 =>
            next_state <= multiplication_with_reduction_special_prime_3_5;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_6;
            end if;
        when multiplication_with_reduction_special_prime_3_6 =>
            next_state <= multiplication_with_reduction_special_prime_3_6;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_7;
            end if;
        when multiplication_with_reduction_special_prime_3_7 =>
            next_state <= multiplication_with_reduction_special_prime_3_7;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_8;
            end if;
        when multiplication_with_reduction_special_prime_3_8 =>
            next_state <= multiplication_with_reduction_special_prime_3_8;
            if(ultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when multiplication_with_reduction_special_prime_3_10 =>
            next_state <= multiplication_with_reduction_special_prime_3_10;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_11;
            end if;
        when multiplication_with_reduction_special_prime_3_11 =>
            next_state <= multiplication_with_reduction_special_prime_3_11;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_12;
            end if;
        when multiplication_with_reduction_special_prime_3_12 =>
            next_state <= multiplication_with_reduction_special_prime_3_12;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_13;
            end if;
        when multiplication_with_reduction_special_prime_3_13 =>
            next_state <= multiplication_with_reduction_special_prime_3_13;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_14;
            end if;
        when multiplication_with_reduction_special_prime_3_14 =>
            next_state <= multiplication_with_reduction_special_prime_3_14;
            if(ultimate_operation = '1') then
                if(operands_size = "011") then
                    next_state <= multiplication_with_reduction_special_prime_3_15;
                else
                    next_state <= multiplication_with_reduction_special_prime_3_27;
                end if;
            end if;
        when multiplication_with_reduction_special_prime_3_15 =>
            next_state <= multiplication_with_reduction_special_prime_3_15;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_16;
            end if;
        when multiplication_with_reduction_special_prime_3_16 =>
            next_state <= multiplication_with_reduction_special_prime_3_16;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_17;
            end if;
        when multiplication_with_reduction_special_prime_3_17 =>
            next_state <= multiplication_with_reduction_special_prime_3_17;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_18;
            end if;
        when multiplication_with_reduction_special_prime_3_18 =>
            next_state <= multiplication_with_reduction_special_prime_3_18;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_19;
            end if;
        when multiplication_with_reduction_special_prime_3_19 =>
            next_state <= multiplication_with_reduction_special_prime_3_19;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_20;
            end if;
        when multiplication_with_reduction_special_prime_3_20 =>
            next_state <= multiplication_with_reduction_special_prime_3_20;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_21;
            end if;
        when multiplication_with_reduction_special_prime_3_21 =>
            next_state <= multiplication_with_reduction_special_prime_3_21;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_22;
            end if;
        when multiplication_with_reduction_special_prime_3_22 =>
            next_state <= multiplication_with_reduction_special_prime_3_22;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_23;
            end if;
        when multiplication_with_reduction_special_prime_3_23 =>
            next_state <= multiplication_with_reduction_special_prime_3_23;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_24;
            end if;
        when multiplication_with_reduction_special_prime_3_24 =>
            next_state <= multiplication_with_reduction_special_prime_3_24;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_25;
            end if;
        when multiplication_with_reduction_special_prime_3_25 =>
            next_state <= multiplication_with_reduction_special_prime_3_25;
            if(ultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when multiplication_with_reduction_special_prime_3_27 =>
            next_state <= multiplication_with_reduction_special_prime_3_27;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_28;
            end if;
        when multiplication_with_reduction_special_prime_3_28 =>
            next_state <= multiplication_with_reduction_special_prime_3_28;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_29;
            end if;
        when multiplication_with_reduction_special_prime_3_29 =>
            next_state <= multiplication_with_reduction_special_prime_3_29;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_30;
            end if;
        when multiplication_with_reduction_special_prime_3_30 =>
            next_state <= multiplication_with_reduction_special_prime_3_30;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_31;
            end if;
        when multiplication_with_reduction_special_prime_3_31 =>
            next_state <= multiplication_with_reduction_special_prime_3_31;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_32;
            end if;
        when multiplication_with_reduction_special_prime_3_32 =>
            next_state <= multiplication_with_reduction_special_prime_3_32;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_33;
            end if;
        when multiplication_with_reduction_special_prime_3_33 =>
            next_state <= multiplication_with_reduction_special_prime_3_33;
            if(ultimate_operation = '1') then
                if(operands_size = "100") then
                    next_state <= multiplication_with_reduction_special_prime_3_34;
                else
                    next_state <= multiplication_with_reduction_special_prime_3_54;
                end if;
            end if;
        when multiplication_with_reduction_special_prime_3_34 =>
            next_state <= multiplication_with_reduction_special_prime_3_34;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_35;
            end if;
        when multiplication_with_reduction_special_prime_3_35 =>
            next_state <= multiplication_with_reduction_special_prime_3_35;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_36;
            end if;
        when multiplication_with_reduction_special_prime_3_36 =>
            next_state <= multiplication_with_reduction_special_prime_3_36;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_37;
            end if;
        when multiplication_with_reduction_special_prime_3_37 =>
            next_state <= multiplication_with_reduction_special_prime_3_37;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_38;
            end if;
        when multiplication_with_reduction_special_prime_3_38 =>
            next_state <= multiplication_with_reduction_special_prime_3_38;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_39;
            end if;
        when multiplication_with_reduction_special_prime_3_39 =>
            next_state <= multiplication_with_reduction_special_prime_3_39;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_40;
            end if;
        when multiplication_with_reduction_special_prime_3_40 =>
            next_state <= multiplication_with_reduction_special_prime_3_40;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_41;
            end if;
        when multiplication_with_reduction_special_prime_3_41 =>
            next_state <= multiplication_with_reduction_special_prime_3_41;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_42;
            end if;
        when multiplication_with_reduction_special_prime_3_42 =>
            next_state <= multiplication_with_reduction_special_prime_3_42;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_43;
            end if;
        when multiplication_with_reduction_special_prime_3_43 =>
            next_state <= multiplication_with_reduction_special_prime_3_43;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_44;
            end if;
        when multiplication_with_reduction_special_prime_3_44 =>
            next_state <= multiplication_with_reduction_special_prime_3_44;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_45;
            end if;
        when multiplication_with_reduction_special_prime_3_45 =>
            next_state <= multiplication_with_reduction_special_prime_3_45;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_46;
            end if;
        when multiplication_with_reduction_special_prime_3_46 =>
            next_state <= multiplication_with_reduction_special_prime_3_46;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_47;
            end if;
        when multiplication_with_reduction_special_prime_3_47 =>
            next_state <= multiplication_with_reduction_special_prime_3_47;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_48;
            end if;
        when multiplication_with_reduction_special_prime_3_48 =>
            next_state <= multiplication_with_reduction_special_prime_3_48;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_49;
            end if;
        when multiplication_with_reduction_special_prime_3_49 =>
            next_state <= multiplication_with_reduction_special_prime_3_49;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_50;
            end if;
        when multiplication_with_reduction_special_prime_3_50 =>
            next_state <= multiplication_with_reduction_special_prime_3_50;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_51;
            end if;
        when multiplication_with_reduction_special_prime_3_51 =>
            next_state <= multiplication_with_reduction_special_prime_3_51;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_52;
            end if;
        when multiplication_with_reduction_special_prime_3_52 =>
            next_state <= multiplication_with_reduction_special_prime_3_52;
            if(ultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when multiplication_with_reduction_special_prime_3_54 =>
            next_state <= multiplication_with_reduction_special_prime_3_54;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_55;
            end if;
        when multiplication_with_reduction_special_prime_3_55 =>
            next_state <= multiplication_with_reduction_special_prime_3_55;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_56;
            end if;
        when multiplication_with_reduction_special_prime_3_56 =>
            next_state <= multiplication_with_reduction_special_prime_3_56;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_57;
            end if;
        when multiplication_with_reduction_special_prime_3_57 =>
            next_state <= multiplication_with_reduction_special_prime_3_57;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_58;
            end if;
        when multiplication_with_reduction_special_prime_3_58 =>
            next_state <= multiplication_with_reduction_special_prime_3_58;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_59;
            end if;
        when multiplication_with_reduction_special_prime_3_59 =>
            next_state <= multiplication_with_reduction_special_prime_3_59;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_60;
            end if;
        when multiplication_with_reduction_special_prime_3_60 =>
            next_state <= multiplication_with_reduction_special_prime_3_60;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_61;
            end if;
        when multiplication_with_reduction_special_prime_3_61 =>
            next_state <= multiplication_with_reduction_special_prime_3_61;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_62;
            end if;
        when multiplication_with_reduction_special_prime_3_62 =>
            next_state <= multiplication_with_reduction_special_prime_3_62;
            if(ultimate_operation = '1') then
                if(operands_size = "101") then
                    next_state <= multiplication_with_reduction_special_prime_3_63;
                else
                    next_state <= multiplication_with_reduction_special_prime_3_93;
                end if;
            end if;
        when multiplication_with_reduction_special_prime_3_63 =>
            next_state <= multiplication_with_reduction_special_prime_3_63;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_64;
            end if;
        when multiplication_with_reduction_special_prime_3_64 =>
            next_state <= multiplication_with_reduction_special_prime_3_64;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_65;
            end if;
        when multiplication_with_reduction_special_prime_3_65 =>
            next_state <= multiplication_with_reduction_special_prime_3_65;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_66;
            end if;
        when multiplication_with_reduction_special_prime_3_66 =>
            next_state <= multiplication_with_reduction_special_prime_3_66;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_67;
            end if;
        when multiplication_with_reduction_special_prime_3_67 =>
            next_state <= multiplication_with_reduction_special_prime_3_67;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_68;
            end if;
        when multiplication_with_reduction_special_prime_3_68 =>
            next_state <= multiplication_with_reduction_special_prime_3_68;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_69;
            end if;
        when multiplication_with_reduction_special_prime_3_69 =>
            next_state <= multiplication_with_reduction_special_prime_3_69;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_70;
            end if;
        when multiplication_with_reduction_special_prime_3_70 =>
            next_state <= multiplication_with_reduction_special_prime_3_70;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_71;
            end if;
        when multiplication_with_reduction_special_prime_3_71 =>
            next_state <= multiplication_with_reduction_special_prime_3_71;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_72;
            end if;
        when multiplication_with_reduction_special_prime_3_72 =>
            next_state <= multiplication_with_reduction_special_prime_3_72;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_73;
            end if;
        when multiplication_with_reduction_special_prime_3_73 =>
            next_state <= multiplication_with_reduction_special_prime_3_73;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_74;
            end if;
        when multiplication_with_reduction_special_prime_3_74 =>
            next_state <= multiplication_with_reduction_special_prime_3_74;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_75;
            end if;
        when multiplication_with_reduction_special_prime_3_75 =>
            next_state <= multiplication_with_reduction_special_prime_3_75;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_76;
            end if;
        when multiplication_with_reduction_special_prime_3_76 =>
            next_state <= multiplication_with_reduction_special_prime_3_76;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_77;
            end if;
        when multiplication_with_reduction_special_prime_3_77 =>
            next_state <= multiplication_with_reduction_special_prime_3_77;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_78;
            end if;
        when multiplication_with_reduction_special_prime_3_78 =>
            next_state <= multiplication_with_reduction_special_prime_3_78;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_79;
            end if;
        when multiplication_with_reduction_special_prime_3_79 =>
            next_state <= multiplication_with_reduction_special_prime_3_79;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_80;
            end if;
        when multiplication_with_reduction_special_prime_3_80 =>
            next_state <= multiplication_with_reduction_special_prime_3_80;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_81;
            end if;
        when multiplication_with_reduction_special_prime_3_81 =>
            next_state <= multiplication_with_reduction_special_prime_3_81;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_82;
            end if;
        when multiplication_with_reduction_special_prime_3_82 =>
            next_state <= multiplication_with_reduction_special_prime_3_82;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_83;
            end if;
        when multiplication_with_reduction_special_prime_3_83 =>
            next_state <= multiplication_with_reduction_special_prime_3_83;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_84;
            end if;
        when multiplication_with_reduction_special_prime_3_84 =>
            next_state <= multiplication_with_reduction_special_prime_3_84;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_85;
            end if;
        when multiplication_with_reduction_special_prime_3_85 =>
            next_state <= multiplication_with_reduction_special_prime_3_85;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_86;
            end if;
        when multiplication_with_reduction_special_prime_3_86 =>
            next_state <= multiplication_with_reduction_special_prime_3_86;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_87;
            end if;
        when multiplication_with_reduction_special_prime_3_87 =>
            next_state <= multiplication_with_reduction_special_prime_3_87;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_88;
            end if;
        when multiplication_with_reduction_special_prime_3_88 =>
            next_state <= multiplication_with_reduction_special_prime_3_88;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_89;
            end if;
        when multiplication_with_reduction_special_prime_3_89 =>
            next_state <= multiplication_with_reduction_special_prime_3_89;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_90;
            end if;
        when multiplication_with_reduction_special_prime_3_90 =>
            next_state <= multiplication_with_reduction_special_prime_3_90;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_91;
            end if;
        when multiplication_with_reduction_special_prime_3_91 =>
            next_state <= multiplication_with_reduction_special_prime_3_91;
            if(ultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when multiplication_with_reduction_special_prime_3_93 =>
            next_state <= multiplication_with_reduction_special_prime_3_93;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_94;
            end if;
        when multiplication_with_reduction_special_prime_3_94 =>
            next_state <= multiplication_with_reduction_special_prime_3_94;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_95;
            end if;
        when multiplication_with_reduction_special_prime_3_95 =>
            next_state <= multiplication_with_reduction_special_prime_3_95;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_96;
            end if;
        when multiplication_with_reduction_special_prime_3_96 =>
            next_state <= multiplication_with_reduction_special_prime_3_96;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_97;
            end if;
        when multiplication_with_reduction_special_prime_3_97 =>
            next_state <= multiplication_with_reduction_special_prime_3_97;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_98;
            end if;
        when multiplication_with_reduction_special_prime_3_98 =>
            next_state <= multiplication_with_reduction_special_prime_3_98;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_99;
            end if;
        when multiplication_with_reduction_special_prime_3_99 =>
            next_state <= multiplication_with_reduction_special_prime_3_99;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_100;
            end if;
        when multiplication_with_reduction_special_prime_3_100 =>
            next_state <= multiplication_with_reduction_special_prime_3_100;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_101;
            end if;
        when multiplication_with_reduction_special_prime_3_101 =>
            next_state <= multiplication_with_reduction_special_prime_3_101;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_102;
            end if;
        when multiplication_with_reduction_special_prime_3_102 =>
            next_state <= multiplication_with_reduction_special_prime_3_102;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_103;
            end if;
        when multiplication_with_reduction_special_prime_3_103 => 
            next_state <= multiplication_with_reduction_special_prime_3_103;
            if(ultimate_operation = '1') then
                if(operands_size = "110") then
                    next_state <= multiplication_with_reduction_special_prime_3_104;
                else
                    next_state <= multiplication_with_reduction_special_prime_3_146;
                end if;
            end if;
        when multiplication_with_reduction_special_prime_3_104 => 
            next_state <= multiplication_with_reduction_special_prime_3_104;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_105;
            end if;
        when multiplication_with_reduction_special_prime_3_105 => 
            next_state <= multiplication_with_reduction_special_prime_3_105;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_106;
            end if;
        when multiplication_with_reduction_special_prime_3_106 => 
            next_state <= multiplication_with_reduction_special_prime_3_106;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_107;
            end if;
        when multiplication_with_reduction_special_prime_3_107 => 
            next_state <= multiplication_with_reduction_special_prime_3_107;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_108;
            end if;
        when multiplication_with_reduction_special_prime_3_108 => 
            next_state <= multiplication_with_reduction_special_prime_3_108;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_109;
            end if;
        when multiplication_with_reduction_special_prime_3_109 => 
            next_state <= multiplication_with_reduction_special_prime_3_109;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_110;
            end if;
        when multiplication_with_reduction_special_prime_3_110 => 
            next_state <= multiplication_with_reduction_special_prime_3_110;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_111;
            end if;
        when multiplication_with_reduction_special_prime_3_111 => 
            next_state <= multiplication_with_reduction_special_prime_3_111;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_112;
            end if;
        when multiplication_with_reduction_special_prime_3_112 => 
            next_state <= multiplication_with_reduction_special_prime_3_112;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_113;
            end if;
        when multiplication_with_reduction_special_prime_3_113 => 
            next_state <= multiplication_with_reduction_special_prime_3_113;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_114;
            end if;
        when multiplication_with_reduction_special_prime_3_114 => 
            next_state <= multiplication_with_reduction_special_prime_3_114;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_115;
            end if;
        when multiplication_with_reduction_special_prime_3_115 => 
            next_state <= multiplication_with_reduction_special_prime_3_115;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_116;
            end if;
        when multiplication_with_reduction_special_prime_3_116 => 
            next_state <= multiplication_with_reduction_special_prime_3_116;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_117;
            end if;
        when multiplication_with_reduction_special_prime_3_117 => 
            next_state <= multiplication_with_reduction_special_prime_3_117;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_118;
            end if;
        when multiplication_with_reduction_special_prime_3_118 => 
            next_state <= multiplication_with_reduction_special_prime_3_118;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_119;
            end if;
        when multiplication_with_reduction_special_prime_3_119 => 
            next_state <= multiplication_with_reduction_special_prime_3_119;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_120;
            end if;
        when multiplication_with_reduction_special_prime_3_120 => 
            next_state <= multiplication_with_reduction_special_prime_3_120;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_121;
            end if;
        when multiplication_with_reduction_special_prime_3_121 => 
            next_state <= multiplication_with_reduction_special_prime_3_121;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_122;
            end if;
        when multiplication_with_reduction_special_prime_3_122 => 
            next_state <= multiplication_with_reduction_special_prime_3_122;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_123;
            end if;
        when multiplication_with_reduction_special_prime_3_123 => 
            next_state <= multiplication_with_reduction_special_prime_3_123;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_124;
            end if;
        when multiplication_with_reduction_special_prime_3_124 => 
            next_state <= multiplication_with_reduction_special_prime_3_124;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_125;
            end if;
        when multiplication_with_reduction_special_prime_3_125 => 
            next_state <= multiplication_with_reduction_special_prime_3_125;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_126;
            end if;
        when multiplication_with_reduction_special_prime_3_126 => 
            next_state <= multiplication_with_reduction_special_prime_3_126;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_127;
            end if;
        when multiplication_with_reduction_special_prime_3_127 => 
            next_state <= multiplication_with_reduction_special_prime_3_127;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_128;
            end if;
        when multiplication_with_reduction_special_prime_3_128 => 
            next_state <= multiplication_with_reduction_special_prime_3_128;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_129;
            end if;
        when multiplication_with_reduction_special_prime_3_129 => 
            next_state <= multiplication_with_reduction_special_prime_3_129;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_130;
            end if;
        when multiplication_with_reduction_special_prime_3_130 => 
            next_state <= multiplication_with_reduction_special_prime_3_130;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_131;
            end if;
        when multiplication_with_reduction_special_prime_3_131 => 
            next_state <= multiplication_with_reduction_special_prime_3_131;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_132;
            end if;
        when multiplication_with_reduction_special_prime_3_132 => 
            next_state <= multiplication_with_reduction_special_prime_3_132;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_133;
            end if;
        when multiplication_with_reduction_special_prime_3_133 => 
            next_state <= multiplication_with_reduction_special_prime_3_133;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_134;
            end if;
        when multiplication_with_reduction_special_prime_3_134 => 
            next_state <= multiplication_with_reduction_special_prime_3_134;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_135;
            end if;
        when multiplication_with_reduction_special_prime_3_135 => 
            next_state <= multiplication_with_reduction_special_prime_3_135;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_136;
            end if;
        when multiplication_with_reduction_special_prime_3_136 => 
            next_state <= multiplication_with_reduction_special_prime_3_136;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_137;
            end if;
        when multiplication_with_reduction_special_prime_3_137 => 
            next_state <= multiplication_with_reduction_special_prime_3_137;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_138;
            end if;
        when multiplication_with_reduction_special_prime_3_138 => 
            next_state <= multiplication_with_reduction_special_prime_3_138;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_139;
            end if;
        when multiplication_with_reduction_special_prime_3_139 => 
            next_state <= multiplication_with_reduction_special_prime_3_139;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_140;
            end if;
        when multiplication_with_reduction_special_prime_3_140 => 
            next_state <= multiplication_with_reduction_special_prime_3_140;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_141;
            end if;
        when multiplication_with_reduction_special_prime_3_141 => 
            next_state <= multiplication_with_reduction_special_prime_3_141;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_142;
            end if;
        when multiplication_with_reduction_special_prime_3_142 => 
            next_state <= multiplication_with_reduction_special_prime_3_142;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_143;
            end if;
        when multiplication_with_reduction_special_prime_3_143 => 
            next_state <= multiplication_with_reduction_special_prime_3_143;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_144;
            end if;
        when multiplication_with_reduction_special_prime_3_144 => 
            next_state <= multiplication_with_reduction_special_prime_3_144;
            if(ultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when multiplication_with_reduction_special_prime_3_146 => 
            next_state <= multiplication_with_reduction_special_prime_3_146;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_147;
            end if;
        when multiplication_with_reduction_special_prime_3_147 => 
            next_state <= multiplication_with_reduction_special_prime_3_147;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_148;
            end if;
        when multiplication_with_reduction_special_prime_3_148 => 
            next_state <= multiplication_with_reduction_special_prime_3_148;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_149;
            end if;
        when multiplication_with_reduction_special_prime_3_149 => 
            next_state <= multiplication_with_reduction_special_prime_3_149;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_150;
            end if;
        when multiplication_with_reduction_special_prime_3_150 => 
            next_state <= multiplication_with_reduction_special_prime_3_150;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_151;
            end if;
        when multiplication_with_reduction_special_prime_3_151 => 
            next_state <= multiplication_with_reduction_special_prime_3_151;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_152;
            end if;
        when multiplication_with_reduction_special_prime_3_152 => 
            next_state <= multiplication_with_reduction_special_prime_3_152;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_153;
            end if;
        when multiplication_with_reduction_special_prime_3_153 => 
            next_state <= multiplication_with_reduction_special_prime_3_153;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_154;
            end if;
        when multiplication_with_reduction_special_prime_3_154 => 
            next_state <= multiplication_with_reduction_special_prime_3_154;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_155;
            end if;
        when multiplication_with_reduction_special_prime_3_155 => 
            next_state <= multiplication_with_reduction_special_prime_3_155;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_156;
            end if;
        when multiplication_with_reduction_special_prime_3_156 => 
            next_state <= multiplication_with_reduction_special_prime_3_156;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_157;
            end if;
        when multiplication_with_reduction_special_prime_3_157 => 
            next_state <= multiplication_with_reduction_special_prime_3_157;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_158;
            end if;
        when multiplication_with_reduction_special_prime_3_158 => 
            next_state <= multiplication_with_reduction_special_prime_3_158;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_159;
            end if;
        when multiplication_with_reduction_special_prime_3_159 => 
            next_state <= multiplication_with_reduction_special_prime_3_159;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_160;
            end if;
        when multiplication_with_reduction_special_prime_3_160 => 
            next_state <= multiplication_with_reduction_special_prime_3_160;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_161;
            end if;
        when multiplication_with_reduction_special_prime_3_161 => 
            next_state <= multiplication_with_reduction_special_prime_3_161;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_162;
            end if;
        when multiplication_with_reduction_special_prime_3_162 => 
            next_state <= multiplication_with_reduction_special_prime_3_162;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_163;
            end if;
        when multiplication_with_reduction_special_prime_3_163 => 
            next_state <= multiplication_with_reduction_special_prime_3_163;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_164;
            end if;
        when multiplication_with_reduction_special_prime_3_164 => 
            next_state <= multiplication_with_reduction_special_prime_3_164;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_165;
            end if;
        when multiplication_with_reduction_special_prime_3_165 => 
            next_state <= multiplication_with_reduction_special_prime_3_165;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_166;
            end if;
        when multiplication_with_reduction_special_prime_3_166 => 
            next_state <= multiplication_with_reduction_special_prime_3_166;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_167;
            end if;
        when multiplication_with_reduction_special_prime_3_167 => 
            next_state <= multiplication_with_reduction_special_prime_3_167;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_168;
            end if;
        when multiplication_with_reduction_special_prime_3_168 => 
            next_state <= multiplication_with_reduction_special_prime_3_168;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_169;
            end if;
        when multiplication_with_reduction_special_prime_3_169 => 
            next_state <= multiplication_with_reduction_special_prime_3_169;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_170;
            end if;
        when multiplication_with_reduction_special_prime_3_170 => 
            next_state <= multiplication_with_reduction_special_prime_3_170;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_171;
            end if;
        when multiplication_with_reduction_special_prime_3_171 => 
            next_state <= multiplication_with_reduction_special_prime_3_171;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_172;
            end if;
        when multiplication_with_reduction_special_prime_3_172 => 
            next_state <= multiplication_with_reduction_special_prime_3_172;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_173;
            end if;
        when multiplication_with_reduction_special_prime_3_173 => 
            next_state <= multiplication_with_reduction_special_prime_3_173;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_174;
            end if;
        when multiplication_with_reduction_special_prime_3_174 => 
            next_state <= multiplication_with_reduction_special_prime_3_174;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_175;
            end if;
        when multiplication_with_reduction_special_prime_3_175 => 
            next_state <= multiplication_with_reduction_special_prime_3_175;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_176;
            end if;
        when multiplication_with_reduction_special_prime_3_176 => 
            next_state <= multiplication_with_reduction_special_prime_3_176;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_177;
            end if;
        when multiplication_with_reduction_special_prime_3_177 => 
            next_state <= multiplication_with_reduction_special_prime_3_177;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_178;
            end if;
        when multiplication_with_reduction_special_prime_3_178 => 
            next_state <= multiplication_with_reduction_special_prime_3_178;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_179;
            end if;
        when multiplication_with_reduction_special_prime_3_179 => 
            next_state <= multiplication_with_reduction_special_prime_3_179;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_180;
            end if;
        when multiplication_with_reduction_special_prime_3_180 => 
            next_state <= multiplication_with_reduction_special_prime_3_180;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_181;
            end if;
        when multiplication_with_reduction_special_prime_3_181 => 
            next_state <= multiplication_with_reduction_special_prime_3_181;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_182;
            end if;
        when multiplication_with_reduction_special_prime_3_182 => 
            next_state <= multiplication_with_reduction_special_prime_3_182;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_183;
            end if;
        when multiplication_with_reduction_special_prime_3_183 => 
            next_state <= multiplication_with_reduction_special_prime_3_183;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_184;
            end if;
        when multiplication_with_reduction_special_prime_3_184 => 
            next_state <= multiplication_with_reduction_special_prime_3_184;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_185;
            end if;
        when multiplication_with_reduction_special_prime_3_185 => 
            next_state <= multiplication_with_reduction_special_prime_3_185;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_186;
            end if;
        when multiplication_with_reduction_special_prime_3_186 => 
            next_state <= multiplication_with_reduction_special_prime_3_186;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_187;
            end if;
        when multiplication_with_reduction_special_prime_3_187 => 
            next_state <= multiplication_with_reduction_special_prime_3_187;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_188;
            end if;
        when multiplication_with_reduction_special_prime_3_188 => 
            next_state <= multiplication_with_reduction_special_prime_3_188;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_189;
            end if;
        when multiplication_with_reduction_special_prime_3_189 => 
            next_state <= multiplication_with_reduction_special_prime_3_189;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_190;
            end if;
        when multiplication_with_reduction_special_prime_3_190 => 
            next_state <= multiplication_with_reduction_special_prime_3_190;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_191;
            end if;
        when multiplication_with_reduction_special_prime_3_191 => 
            next_state <= multiplication_with_reduction_special_prime_3_191;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_192;
            end if;
        when multiplication_with_reduction_special_prime_3_192 => 
            next_state <= multiplication_with_reduction_special_prime_3_192;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_193;
            end if;
        when multiplication_with_reduction_special_prime_3_193 => 
            next_state <= multiplication_with_reduction_special_prime_3_193;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_194;
            end if;
        when multiplication_with_reduction_special_prime_3_194 => 
            next_state <= multiplication_with_reduction_special_prime_3_194;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_195;
            end if;
        when multiplication_with_reduction_special_prime_3_195 => 
            next_state <= multiplication_with_reduction_special_prime_3_195;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_196;
            end if;
        when multiplication_with_reduction_special_prime_3_196 => 
            next_state <= multiplication_with_reduction_special_prime_3_196;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_197;
            end if;
        when multiplication_with_reduction_special_prime_3_197 => 
            next_state <= multiplication_with_reduction_special_prime_3_197;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_198;
            end if;
        when multiplication_with_reduction_special_prime_3_198 => 
            next_state <= multiplication_with_reduction_special_prime_3_198;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_199;
            end if;
        when multiplication_with_reduction_special_prime_3_199 => 
            next_state <= multiplication_with_reduction_special_prime_3_199;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_200;
            end if;
        when multiplication_with_reduction_special_prime_3_200 => 
            next_state <= multiplication_with_reduction_special_prime_3_200;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_201;
            end if;
        when multiplication_with_reduction_special_prime_3_201 => 
            next_state <= multiplication_with_reduction_special_prime_3_201;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_202;
            end if;
        when multiplication_with_reduction_special_prime_3_202 => 
            next_state <= multiplication_with_reduction_special_prime_3_202;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_203;
            end if;
        when multiplication_with_reduction_special_prime_3_203 => 
            next_state <= multiplication_with_reduction_special_prime_3_203;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_204;
            end if;
        when multiplication_with_reduction_special_prime_3_204 => 
            next_state <= multiplication_with_reduction_special_prime_3_204;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_205;
            end if;
        when multiplication_with_reduction_special_prime_3_205 => 
            next_state <= multiplication_with_reduction_special_prime_3_205;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_206;
            end if;
        when multiplication_with_reduction_special_prime_3_206 => 
            next_state <= multiplication_with_reduction_special_prime_3_206;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_207;
            end if;
        when multiplication_with_reduction_special_prime_3_207 => 
            next_state <= multiplication_with_reduction_special_prime_3_207;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_208;
            end if;
        when multiplication_with_reduction_special_prime_3_208 => 
            next_state <= multiplication_with_reduction_special_prime_3_208;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_209;
            end if;
        when multiplication_with_reduction_special_prime_3_209 => 
            next_state <= multiplication_with_reduction_special_prime_3_209;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_210;
            end if;
        when multiplication_with_reduction_special_prime_3_210 => 
            next_state <= multiplication_with_reduction_special_prime_3_210;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_211;
            end if;
        when multiplication_with_reduction_special_prime_3_211 => 
            next_state <= multiplication_with_reduction_special_prime_3_211;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_212;
            end if;
        when multiplication_with_reduction_special_prime_3_212 => 
            next_state <= multiplication_with_reduction_special_prime_3_212;
            if(ultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_3_213;
            end if;
        when multiplication_with_reduction_special_prime_3_213 => 
            next_state <= multiplication_with_reduction_special_prime_3_213;
            if(ultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when square_with_reduction_0 => 
            next_state <= square_with_reduction_0;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_1;
            end if;
        when square_with_reduction_1 => 
            next_state <= square_with_reduction_1;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_2;
            end if;
        when square_with_reduction_2 => 
            next_state <= square_with_reduction_2;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_3;
            end if;
        when square_with_reduction_3 => 
            next_state <= square_with_reduction_3;
            if(ultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when square_with_reduction_5 => 
            next_state <= square_with_reduction_5;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_6;
            end if;
        when square_with_reduction_6 => 
            next_state <= square_with_reduction_6;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_7;
            end if;
        when square_with_reduction_7 => 
            next_state <= square_with_reduction_7;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_8;
            end if;
        when square_with_reduction_8 => 
            next_state <= square_with_reduction_8;
            if(ultimate_operation = '1') then
                if(operands_size = "001") then
                    next_state <= square_with_reduction_9;
                else
                    next_state <= square_with_reduction_15;
                end if;
            end if;
        when square_with_reduction_9 => 
            next_state <= square_with_reduction_9;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_10;
            end if;
        when square_with_reduction_10 => 
            next_state <= square_with_reduction_10;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_11;
            end if;
        when square_with_reduction_11 => 
            next_state <= square_with_reduction_11;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_12;
            end if;
        when square_with_reduction_12 => 
            next_state <= square_with_reduction_12;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_13;
            end if;
        when square_with_reduction_13 => 
            next_state <= square_with_reduction_13;
            if(ultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when square_with_reduction_15 => 
            next_state <= square_with_reduction_15;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_16;
            end if;
        when square_with_reduction_16 => 
            next_state <= square_with_reduction_16;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_17;
            end if;
        when square_with_reduction_17 => 
            next_state <= square_with_reduction_17;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_18;
            end if;
        when square_with_reduction_18 => 
            next_state <= square_with_reduction_18;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_19;
            end if;
        when square_with_reduction_19 => 
            next_state <= square_with_reduction_19;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_20;
            end if;
        when square_with_reduction_20 => 
            next_state <= square_with_reduction_20;
            if(ultimate_operation = '1') then
                if(operands_size = "010") then
                    next_state <= square_with_reduction_21;
                else
                    next_state <= square_with_reduction_30;
                end if;
            end if;
        when square_with_reduction_21 => 
            next_state <= square_with_reduction_21;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_22;
            end if;
        when square_with_reduction_22 => 
            next_state <= square_with_reduction_22;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_23;
            end if;
        when square_with_reduction_23 => 
            next_state <= square_with_reduction_23;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_24;
            end if;
        when square_with_reduction_24 => 
            next_state <= square_with_reduction_24;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_25;
            end if;
        when square_with_reduction_25 => 
            next_state <= square_with_reduction_25;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_26;
            end if;
        when square_with_reduction_26 => 
            next_state <= square_with_reduction_26;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_27;
            end if;
        when square_with_reduction_27 => 
            next_state <= square_with_reduction_27;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_28;
            end if;
        when square_with_reduction_28 => 
            next_state <= square_with_reduction_28;
            if(ultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when square_with_reduction_30 => 
            next_state <= square_with_reduction_30;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_31;
            end if;
        when square_with_reduction_31 => 
            next_state <= square_with_reduction_31;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_32;
            end if;
        when square_with_reduction_32 => 
            next_state <= square_with_reduction_32;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_33;
            end if;
        when square_with_reduction_33 => 
            next_state <= square_with_reduction_33;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_34;
            end if;
        when square_with_reduction_34 => 
            next_state <= square_with_reduction_34;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_35;
            end if;
        when square_with_reduction_35 => 
            next_state <= square_with_reduction_35;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_36;
            end if;
        when square_with_reduction_36 => 
            next_state <= square_with_reduction_36;
            if(ultimate_operation = '1') then
                if(operands_size = "011") then
                    next_state <= square_with_reduction_37;
                else
                    next_state <= square_with_reduction_51;
                end if;
            end if;
        when square_with_reduction_37 => 
            next_state <= square_with_reduction_37;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_38;
            end if;
        when square_with_reduction_38 => 
            next_state <= square_with_reduction_38;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_39;
            end if;
        when square_with_reduction_39 => 
            next_state <= square_with_reduction_39;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_40;
            end if;
        when square_with_reduction_40 => 
            next_state <= square_with_reduction_40;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_41;
            end if;
        when square_with_reduction_41 => 
            next_state <= square_with_reduction_41;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_42;
            end if;
        when square_with_reduction_42 => 
            next_state <= square_with_reduction_42;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_43;
            end if;
        when square_with_reduction_43 => 
            next_state <= square_with_reduction_43;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_44;
            end if;
        when square_with_reduction_44 => 
            next_state <= square_with_reduction_44;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_45;
            end if;
        when square_with_reduction_45 => 
            next_state <= square_with_reduction_45;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_46;
            end if;
        when square_with_reduction_46 => 
            next_state <= square_with_reduction_46;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_47;
            end if;
        when square_with_reduction_47 => 
            next_state <= square_with_reduction_47;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_48;
            end if;
        when square_with_reduction_48 => 
            next_state <= square_with_reduction_48;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_49;
            end if;
        when square_with_reduction_49 => 
            next_state <= square_with_reduction_49;
            if(ultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when square_with_reduction_51 => 
            next_state <= square_with_reduction_51;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_52;
            end if;
        when square_with_reduction_52 => 
            next_state <= square_with_reduction_52;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_53;
            end if;
        when square_with_reduction_53 => 
            next_state <= square_with_reduction_53;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_54;
            end if;
        when square_with_reduction_54 => 
            next_state <= square_with_reduction_54;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_55;
            end if;
        when square_with_reduction_55 => 
            next_state <= square_with_reduction_55;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_56;
            end if;
        when square_with_reduction_56 => 
            next_state <= square_with_reduction_56;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_57;
            end if;
        when square_with_reduction_57 => 
            next_state <= square_with_reduction_57;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_58;
            end if;
        when square_with_reduction_58 => 
            next_state <= square_with_reduction_58;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_59;
            end if;
        when square_with_reduction_59 => 
            next_state <= square_with_reduction_59;
            if(ultimate_operation = '1') then
                if(operands_size = "100") then
                    next_state <= square_with_reduction_60;
                else
                    next_state <= square_with_reduction_80;
                end if;
            end if;
        when square_with_reduction_60 => 
            next_state <= square_with_reduction_60;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_61;
            end if;
        when square_with_reduction_61 => 
            next_state <= square_with_reduction_61;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_62;
            end if;
        when square_with_reduction_62 => 
            next_state <= square_with_reduction_62;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_63;
            end if;
        when square_with_reduction_63 => 
            next_state <= square_with_reduction_63;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_64;
            end if;
        when square_with_reduction_64 => 
            next_state <= square_with_reduction_64;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_65;
            end if;
        when square_with_reduction_65 => 
            next_state <= square_with_reduction_65;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_66;
            end if;
        when square_with_reduction_66 => 
            next_state <= square_with_reduction_66;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_67;
            end if;
        when square_with_reduction_67 => 
            next_state <= square_with_reduction_67;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_68;
            end if;
        when square_with_reduction_68 => 
            next_state <= square_with_reduction_68;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_69;
            end if;
        when square_with_reduction_69 => 
            next_state <= square_with_reduction_69;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_70;
            end if;
        when square_with_reduction_70 => 
            next_state <= square_with_reduction_70;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_71;
            end if;
        when square_with_reduction_71 => 
            next_state <= square_with_reduction_71;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_72;
            end if;
        when square_with_reduction_72 => 
            next_state <= square_with_reduction_72;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_73;
            end if;
        when square_with_reduction_73 => 
            next_state <= square_with_reduction_73;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_74;
            end if;
        when square_with_reduction_74 => 
            next_state <= square_with_reduction_74;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_75;
            end if;
        when square_with_reduction_75 => 
            next_state <= square_with_reduction_75;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_76;
            end if;
        when square_with_reduction_76 => 
            next_state <= square_with_reduction_76;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_77;
            end if;
        when square_with_reduction_77 => 
            next_state <= square_with_reduction_77;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_78;
            end if;
        when square_with_reduction_78 => 
            next_state <= square_with_reduction_78;
            if(ultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when square_with_reduction_80 => 
            next_state <= square_with_reduction_80;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_81;
            end if;
        when square_with_reduction_81 => 
            next_state <= square_with_reduction_81;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_82;
            end if;
        when square_with_reduction_82 => 
            next_state <= square_with_reduction_82;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_83;
            end if;
        when square_with_reduction_83 => 
            next_state <= square_with_reduction_83;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_84;
            end if;
        when square_with_reduction_84 => 
            next_state <= square_with_reduction_84;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_85;
            end if;
        when square_with_reduction_85 => 
            next_state <= square_with_reduction_85;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_86;
            end if;
        when square_with_reduction_86 => 
            next_state <= square_with_reduction_86;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_87;
            end if;
        when square_with_reduction_87 => 
            next_state <= square_with_reduction_87;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_88;
            end if;
        when square_with_reduction_88 => 
            next_state <= square_with_reduction_88;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_89;
            end if;
        when square_with_reduction_89 => 
            next_state <= square_with_reduction_89;
            if(ultimate_operation = '1') then
                if(operands_size = "101") then
                    next_state <= square_with_reduction_90;
                else
                    next_state <= square_with_reduction_118;
                end if;
            end if;
        when square_with_reduction_90 => 
            next_state <= square_with_reduction_90;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_91;
            end if;
        when square_with_reduction_91 => 
            next_state <= square_with_reduction_91;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_92;
            end if;
        when square_with_reduction_92 => 
            next_state <= square_with_reduction_92;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_93;
            end if;
        when square_with_reduction_93 => 
            next_state <= square_with_reduction_93;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_94;
            end if;
        when square_with_reduction_94 => 
            next_state <= square_with_reduction_94;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_95;
            end if;
        when square_with_reduction_95 => 
            next_state <= square_with_reduction_95;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_96;
            end if;
        when square_with_reduction_96 => 
            next_state <= square_with_reduction_96;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_97;
            end if;
        when square_with_reduction_97 => 
            next_state <= square_with_reduction_97;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_98;
            end if;
        when square_with_reduction_98 => 
            next_state <= square_with_reduction_98;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_99;
            end if;
        when square_with_reduction_99 => 
            next_state <= square_with_reduction_99;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_100;
            end if;
        when square_with_reduction_100 => 
            next_state <= square_with_reduction_100;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_101;
            end if;
        when square_with_reduction_101 => 
            next_state <= square_with_reduction_101;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_102;
            end if;
        when square_with_reduction_102 => 
            next_state <= square_with_reduction_102;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_103;
            end if;
        when square_with_reduction_103 => 
            next_state <= square_with_reduction_103;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_104;
            end if;
        when square_with_reduction_104 => 
            next_state <= square_with_reduction_104;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_105;
            end if;
        when square_with_reduction_105 => 
            next_state <= square_with_reduction_105;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_106;
            end if;
        when square_with_reduction_106 => 
            next_state <= square_with_reduction_106;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_107;
            end if;
        when square_with_reduction_107 => 
            next_state <= square_with_reduction_107;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_108;
            end if;
        when square_with_reduction_108 => 
            next_state <= square_with_reduction_108;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_109;
            end if;
        when square_with_reduction_109 => 
            next_state <= square_with_reduction_109;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_110;
            end if;
        when square_with_reduction_110 => 
            next_state <= square_with_reduction_110;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_111;
            end if;
        when square_with_reduction_111 => 
            next_state <= square_with_reduction_111;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_112;
            end if;
        when square_with_reduction_112 => 
            next_state <= square_with_reduction_112;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_113;
            end if;
        when square_with_reduction_113 => 
            next_state <= square_with_reduction_113;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_114;
            end if;
        when square_with_reduction_114 => 
            next_state <= square_with_reduction_114;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_115;
            end if;
        when square_with_reduction_115 => 
            next_state <= square_with_reduction_115;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_116;
            end if;
        when square_with_reduction_116 => 
            next_state <= square_with_reduction_116;
            if(ultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when square_with_reduction_118 => 
            next_state <= square_with_reduction_118;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_119;
            end if;
        when square_with_reduction_119 => 
            next_state <= square_with_reduction_119;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_120;
            end if;
        when square_with_reduction_120 => 
            next_state <= square_with_reduction_120;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_121;
            end if;
        when square_with_reduction_121 => 
            next_state <= square_with_reduction_121;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_122;
            end if;
        when square_with_reduction_122 => 
            next_state <= square_with_reduction_122;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_123;
            end if;
        when square_with_reduction_123 => 
            next_state <= square_with_reduction_123;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_124;
            end if;
        when square_with_reduction_124 => 
            next_state <= square_with_reduction_124;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_125;
            end if;
        when square_with_reduction_125 => 
            next_state <= square_with_reduction_125;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_126;
            end if;
        when square_with_reduction_126 => 
            next_state <= square_with_reduction_126;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_127;
            end if;
        when square_with_reduction_127 => 
            next_state <= square_with_reduction_127;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_128;
            end if;
        when square_with_reduction_128 => 
            next_state <= square_with_reduction_128;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_129;
            end if;
        when square_with_reduction_129 => 
            next_state <= square_with_reduction_129;
            if(ultimate_operation = '1') then
                if(operands_size = "110") then
                    next_state <= square_with_reduction_130;
                else
                    next_state <= square_with_reduction_167;
                end if;
            end if;
        when square_with_reduction_130 => 
            next_state <= square_with_reduction_130;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_131;
            end if;
        when square_with_reduction_131 => 
            next_state <= square_with_reduction_131;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_132;
            end if;
        when square_with_reduction_132 => 
            next_state <= square_with_reduction_132;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_133;
            end if;
        when square_with_reduction_133 => 
            next_state <= square_with_reduction_133;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_134;
            end if;
        when square_with_reduction_134 => 
            next_state <= square_with_reduction_134;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_135;
            end if;
        when square_with_reduction_135 => 
            next_state <= square_with_reduction_135;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_136;
            end if;
        when square_with_reduction_136 => 
            next_state <= square_with_reduction_136;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_137;
            end if;
        when square_with_reduction_137 => 
            next_state <= square_with_reduction_137;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_138;
            end if;
        when square_with_reduction_138 => 
            next_state <= square_with_reduction_138;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_139;
            end if;
        when square_with_reduction_139 => 
            next_state <= square_with_reduction_139;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_140;
            end if;
        when square_with_reduction_140 => 
            next_state <= square_with_reduction_140;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_141;
            end if;
        when square_with_reduction_141 => 
            next_state <= square_with_reduction_141;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_142;
            end if;
        when square_with_reduction_142 => 
            next_state <= square_with_reduction_142;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_143;
            end if;
        when square_with_reduction_143 => 
            next_state <= square_with_reduction_143;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_144;
            end if;
        when square_with_reduction_144 => 
            next_state <= square_with_reduction_144;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_145;
            end if;
        when square_with_reduction_145 => 
            next_state <= square_with_reduction_145;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_146;
            end if;
        when square_with_reduction_146 => 
            next_state <= square_with_reduction_146;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_147;
            end if;
        when square_with_reduction_147 => 
            next_state <= square_with_reduction_147;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_148;
            end if;
        when square_with_reduction_148 => 
            next_state <= square_with_reduction_148;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_149;
            end if;
        when square_with_reduction_149 => 
            next_state <= square_with_reduction_149;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_150;
            end if;
        when square_with_reduction_150 => 
            next_state <= square_with_reduction_150;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_151;
            end if;
        when square_with_reduction_151 => 
            next_state <= square_with_reduction_151;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_152;
            end if;
        when square_with_reduction_152 => 
            next_state <= square_with_reduction_152;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_153;
            end if;
        when square_with_reduction_153 => 
            next_state <= square_with_reduction_153;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_154;
            end if;
        when square_with_reduction_154 => 
            next_state <= square_with_reduction_154;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_155;
            end if;
        when square_with_reduction_155 => 
            next_state <= square_with_reduction_155;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_156;
            end if;
        when square_with_reduction_156 => 
            next_state <= square_with_reduction_156;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_157;
            end if;
        when square_with_reduction_157 => 
            next_state <= square_with_reduction_157;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_158;
            end if;
        when square_with_reduction_158 => 
            next_state <= square_with_reduction_158;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_159;
            end if;
        when square_with_reduction_159 => 
            next_state <= square_with_reduction_159;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_160;
            end if;
        when square_with_reduction_160 => 
            next_state <= square_with_reduction_160;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_161;
            end if;
        when square_with_reduction_161 => 
            next_state <= square_with_reduction_161;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_162;
            end if;
        when square_with_reduction_162 => 
            next_state <= square_with_reduction_162;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_163;
            end if;
        when square_with_reduction_163 => 
            next_state <= square_with_reduction_163;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_164;
            end if;
        when square_with_reduction_164 => 
            next_state <= square_with_reduction_164;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_165;
            end if;
        when square_with_reduction_165 => 
            next_state <= square_with_reduction_165;
            if(ultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when square_with_reduction_167 => 
            next_state <= square_with_reduction_167;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_168;
            end if;
        when square_with_reduction_168 => 
            next_state <= square_with_reduction_168;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_169;
            end if;
        when square_with_reduction_169 => 
            next_state <= square_with_reduction_169;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_170;
            end if;
        when square_with_reduction_170 => 
            next_state <= square_with_reduction_170;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_171;
            end if;
        when square_with_reduction_171 => 
            next_state <= square_with_reduction_171;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_172;
            end if;
        when square_with_reduction_172 => 
            next_state <= square_with_reduction_172;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_173;
            end if;
        when square_with_reduction_173 => 
            next_state <= square_with_reduction_173;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_174;
            end if;
        when square_with_reduction_174 => 
            next_state <= square_with_reduction_174;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_175;
            end if;
        when square_with_reduction_175 => 
            next_state <= square_with_reduction_175;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_176;
            end if;
        when square_with_reduction_176 => 
            next_state <= square_with_reduction_176;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_177;
            end if;
        when square_with_reduction_177 => 
            next_state <= square_with_reduction_177;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_178;
            end if;
        when square_with_reduction_178 => 
            next_state <= square_with_reduction_178;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_179;
            end if;
        when square_with_reduction_179 => 
            next_state <= square_with_reduction_179;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_180;
            end if;
        when square_with_reduction_180 => 
            next_state <= square_with_reduction_180;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_181;
            end if;
        when square_with_reduction_181 => 
            next_state <= square_with_reduction_181;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_182;
            end if;
        when square_with_reduction_182 => 
            next_state <= square_with_reduction_182;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_183;
            end if;
        when square_with_reduction_183 => 
            next_state <= square_with_reduction_183;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_184;
            end if;
        when square_with_reduction_184 => 
            next_state <= square_with_reduction_184;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_185;
            end if;
        when square_with_reduction_185 => 
            next_state <= square_with_reduction_185;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_186;
            end if;
        when square_with_reduction_186 => 
            next_state <= square_with_reduction_186;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_187;
            end if;
        when square_with_reduction_187 => 
            next_state <= square_with_reduction_187;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_188;
            end if;
        when square_with_reduction_188 => 
            next_state <= square_with_reduction_188;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_189;
            end if;
        when square_with_reduction_189 => 
            next_state <= square_with_reduction_189;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_190;
            end if;
        when square_with_reduction_190 => 
            next_state <= square_with_reduction_190;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_191;
            end if;
        when square_with_reduction_191 => 
            next_state <= square_with_reduction_191;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_192;
            end if;
        when square_with_reduction_192 => 
            next_state <= square_with_reduction_192;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_193;
            end if;
        when square_with_reduction_193 => 
            next_state <= square_with_reduction_193;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_194;
            end if;
        when square_with_reduction_194 => 
            next_state <= square_with_reduction_194;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_195;
            end if;
        when square_with_reduction_195 => 
            next_state <= square_with_reduction_195;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_196;
            end if;
        when square_with_reduction_196 => 
            next_state <= square_with_reduction_196;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_197;
            end if;
        when square_with_reduction_197 => 
            next_state <= square_with_reduction_197;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_198;
            end if;
        when square_with_reduction_198 => 
            next_state <= square_with_reduction_198;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_199;
            end if;
        when square_with_reduction_199 => 
            next_state <= square_with_reduction_199;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_200;
            end if;
        when square_with_reduction_200 => 
            next_state <= square_with_reduction_200;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_201;
            end if;
        when square_with_reduction_201 => 
            next_state <= square_with_reduction_201;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_202;
            end if;
        when square_with_reduction_202 => 
            next_state <= square_with_reduction_202;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_203;
            end if;
        when square_with_reduction_203 => 
            next_state <= square_with_reduction_203;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_204;
            end if;
        when square_with_reduction_204 => 
            next_state <= square_with_reduction_204;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_205;
            end if;
        when square_with_reduction_205 => 
            next_state <= square_with_reduction_205;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_206;
            end if;
        when square_with_reduction_206 => 
            next_state <= square_with_reduction_206;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_207;
            end if;
        when square_with_reduction_207 => 
            next_state <= square_with_reduction_207;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_208;
            end if;
        when square_with_reduction_208 => 
            next_state <= square_with_reduction_208;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_209;
            end if;
        when square_with_reduction_209 => 
            next_state <= square_with_reduction_209;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_210;
            end if;
        when square_with_reduction_210 => 
            next_state <= square_with_reduction_210;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_211;
            end if;
        when square_with_reduction_211 => 
            next_state <= square_with_reduction_211;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_212;
            end if;
        when square_with_reduction_212 => 
            next_state <= square_with_reduction_212;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_213;
            end if;
        when square_with_reduction_213 => 
            next_state <= square_with_reduction_213;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_214;
            end if;
        when square_with_reduction_214 => 
            next_state <= square_with_reduction_214;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_215;
            end if;
        when square_with_reduction_215 => 
            next_state <= square_with_reduction_215;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_216;
            end if;
        when square_with_reduction_216 => 
            next_state <= square_with_reduction_216;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_217;
            end if;
        when square_with_reduction_217 => 
            next_state <= square_with_reduction_217;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_218;
            end if;
        when square_with_reduction_218 => 
            next_state <= square_with_reduction_218;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_219;
            end if;
        when square_with_reduction_219 => 
            next_state <= square_with_reduction_219;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_220;
            end if;
        when square_with_reduction_220 => 
            next_state <= square_with_reduction_220;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_221;
            end if;
        when square_with_reduction_221 => 
            next_state <= square_with_reduction_221;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_222;
            end if;
        when square_with_reduction_222 => 
            next_state <= square_with_reduction_222;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_223;
            end if;
        when square_with_reduction_223 => 
            next_state <= square_with_reduction_223;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_224;
            end if;
        when square_with_reduction_224 => 
            next_state <= square_with_reduction_224;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_225;
            end if;
        when square_with_reduction_225 => 
            next_state <= square_with_reduction_225;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_226;
            end if;
        when square_with_reduction_226 => 
            next_state <= square_with_reduction_226;
            if(ultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when square_with_reduction_special_prime_1_0 => 
            next_state <= square_with_reduction_special_prime_1_0;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_1;
            end if;
        when square_with_reduction_special_prime_1_1 => 
            next_state <= square_with_reduction_special_prime_1_1;
            if(ultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when square_with_reduction_special_prime_1_3 => 
            next_state <= square_with_reduction_special_prime_1_3;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_4;
            end if;
        when square_with_reduction_special_prime_1_4 =>
            next_state <= square_with_reduction_special_prime_1_4;
            if(ultimate_operation = '1') then
                if(operands_size = "001") then
                    next_state <= square_with_reduction_special_prime_1_5;
                else
                    next_state <= square_with_reduction_special_prime_1_9;
                end if;
            end if;
        when square_with_reduction_special_prime_1_5 => 
            next_state <= square_with_reduction_special_prime_1_5;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_6;
            end if;
        when square_with_reduction_special_prime_1_6 => 
            next_state <= square_with_reduction_special_prime_1_6;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_7;
            end if;
        when square_with_reduction_special_prime_1_7 => 
            next_state <= square_with_reduction_special_prime_1_7;
            if(ultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when square_with_reduction_special_prime_1_9 => 
            next_state <= square_with_reduction_special_prime_1_9;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_10;
            end if;
        when square_with_reduction_special_prime_1_10 => 
            next_state <= square_with_reduction_special_prime_1_10;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_11;
            end if;
        when square_with_reduction_special_prime_1_11 => 
            next_state <= square_with_reduction_special_prime_1_11;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_12;
            end if;
        when square_with_reduction_special_prime_1_12 => 
            next_state <= square_with_reduction_special_prime_1_12;
            if(ultimate_operation = '1') then
                if(operands_size = "010") then
                    next_state <= square_with_reduction_special_prime_1_13;
                else
                    next_state <= square_with_reduction_special_prime_1_20;
                end if;
            end if;
        when square_with_reduction_special_prime_1_13 => 
            next_state <= square_with_reduction_special_prime_1_13;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_14;
            end if;
        when square_with_reduction_special_prime_1_14 => 
            next_state <= square_with_reduction_special_prime_1_14;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_15;
            end if;
        when square_with_reduction_special_prime_1_15 => 
            next_state <= square_with_reduction_special_prime_1_15;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_16;
            end if;
        when square_with_reduction_special_prime_1_16 => 
            next_state <= square_with_reduction_special_prime_1_16;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_17;
            end if;
        when square_with_reduction_special_prime_1_17 => 
            next_state <= square_with_reduction_special_prime_1_17;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_18;
            end if;
        when square_with_reduction_special_prime_1_18 => 
            next_state <= square_with_reduction_special_prime_1_18;
            if(ultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when square_with_reduction_special_prime_1_20 => 
            next_state <= square_with_reduction_special_prime_1_20;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_21;
            end if;
        when square_with_reduction_special_prime_1_21 => 
            next_state <= square_with_reduction_special_prime_1_21;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_22;
            end if;
        when square_with_reduction_special_prime_1_22 => 
            next_state <= square_with_reduction_special_prime_1_22;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_23;
            end if;
        when square_with_reduction_special_prime_1_23 => 
            next_state <= square_with_reduction_special_prime_1_23;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_24;
            end if;
        when square_with_reduction_special_prime_1_24 => 
            next_state <= square_with_reduction_special_prime_1_24;
            if(ultimate_operation = '1') then
                if(operands_size = "011") then
                    next_state <= square_with_reduction_special_prime_1_25;
                else
                    next_state <= square_with_reduction_special_prime_1_37;
                end if;
            end if;
        when square_with_reduction_special_prime_1_25 => 
            next_state <= square_with_reduction_special_prime_1_25;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_26;
            end if;
        when square_with_reduction_special_prime_1_26 => 
            next_state <= square_with_reduction_special_prime_1_26;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_27;
            end if;
        when square_with_reduction_special_prime_1_27 => 
            next_state <= square_with_reduction_special_prime_1_27;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_28;
            end if;
        when square_with_reduction_special_prime_1_28 => 
            next_state <= square_with_reduction_special_prime_1_28;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_29;
            end if;
        when square_with_reduction_special_prime_1_29 => 
            next_state <= square_with_reduction_special_prime_1_29;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_30;
            end if;
        when square_with_reduction_special_prime_1_30 => 
            next_state <= square_with_reduction_special_prime_1_30;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_31;
            end if;
        when square_with_reduction_special_prime_1_31 => 
            next_state <= square_with_reduction_special_prime_1_31;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_32;
            end if;
        when square_with_reduction_special_prime_1_32 => 
            next_state <= square_with_reduction_special_prime_1_32;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_33;
            end if;
        when square_with_reduction_special_prime_1_33 => 
            next_state <= square_with_reduction_special_prime_1_33;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_34;
            end if;
        when square_with_reduction_special_prime_1_34 => 
            next_state <= square_with_reduction_special_prime_1_34;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_35;
            end if;
        when square_with_reduction_special_prime_1_35 => 
            next_state <= square_with_reduction_special_prime_1_35;
            if(ultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when square_with_reduction_special_prime_1_37 =>
            next_state <= square_with_reduction_special_prime_1_37;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_38;
            end if;
        when square_with_reduction_special_prime_1_38 =>
            next_state <= square_with_reduction_special_prime_1_38;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_39;
            end if;
        when square_with_reduction_special_prime_1_39 =>
            next_state <= square_with_reduction_special_prime_1_39;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_40;
            end if;
        when square_with_reduction_special_prime_1_40 =>
            next_state <= square_with_reduction_special_prime_1_40;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_41;
            end if;
        when square_with_reduction_special_prime_1_41 =>
            next_state <= square_with_reduction_special_prime_1_41;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_42;
            end if;
        when square_with_reduction_special_prime_1_42 =>
            next_state <= square_with_reduction_special_prime_1_42;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_43;
            end if;
        when square_with_reduction_special_prime_1_43 =>
            next_state <= square_with_reduction_special_prime_1_43;
            if(ultimate_operation = '1') then
                if(operands_size = "100") then
                    next_state <= square_with_reduction_special_prime_1_44;
                else
                    next_state <= square_with_reduction_special_prime_1_62;
                end if;
            end if;
        when square_with_reduction_special_prime_1_44 =>
            next_state <= square_with_reduction_special_prime_1_44;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_45;
            end if;
        when square_with_reduction_special_prime_1_45 =>
            next_state <= square_with_reduction_special_prime_1_45;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_46;
            end if;
        when square_with_reduction_special_prime_1_46 =>
            next_state <= square_with_reduction_special_prime_1_46;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_47;
            end if;
        when square_with_reduction_special_prime_1_47 =>
            next_state <= square_with_reduction_special_prime_1_47;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_48;
            end if;
        when square_with_reduction_special_prime_1_48 =>
            next_state <= square_with_reduction_special_prime_1_48;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_49;
            end if;
        when square_with_reduction_special_prime_1_49 =>
            next_state <= square_with_reduction_special_prime_1_49;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_50;
            end if;
        when square_with_reduction_special_prime_1_50 =>
            next_state <= square_with_reduction_special_prime_1_50;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_51;
            end if;
        when square_with_reduction_special_prime_1_51 =>
            next_state <= square_with_reduction_special_prime_1_51;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_52;
            end if;
        when square_with_reduction_special_prime_1_52 =>
            next_state <= square_with_reduction_special_prime_1_52;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_53;
            end if;
        when square_with_reduction_special_prime_1_53 =>
            next_state <= square_with_reduction_special_prime_1_53;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_54;
            end if;
        when square_with_reduction_special_prime_1_54 =>
            next_state <= square_with_reduction_special_prime_1_54;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_55;
            end if;
        when square_with_reduction_special_prime_1_55 =>
            next_state <= square_with_reduction_special_prime_1_55;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_56;
            end if;
        when square_with_reduction_special_prime_1_56 =>
            next_state <= square_with_reduction_special_prime_1_56;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_57;
            end if;
        when square_with_reduction_special_prime_1_57 =>
            next_state <= square_with_reduction_special_prime_1_57;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_58;
            end if;
        when square_with_reduction_special_prime_1_58 =>
            next_state <= square_with_reduction_special_prime_1_58;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_59;
            end if;
        when square_with_reduction_special_prime_1_59 =>
            next_state <= square_with_reduction_special_prime_1_59;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_60;
            end if;
        when square_with_reduction_special_prime_1_60 =>
            next_state <= square_with_reduction_special_prime_1_60;
            if(ultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when square_with_reduction_special_prime_1_62 =>
            next_state <= square_with_reduction_special_prime_1_62;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_63;
            end if;
        when square_with_reduction_special_prime_1_63 =>
            next_state <= square_with_reduction_special_prime_1_63;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_64;
            end if;
        when square_with_reduction_special_prime_1_64 =>
            next_state <= square_with_reduction_special_prime_1_64;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_65;
            end if;
        when square_with_reduction_special_prime_1_65 =>
            next_state <= square_with_reduction_special_prime_1_65;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_66;
            end if;
        when square_with_reduction_special_prime_1_66 =>
            next_state <= square_with_reduction_special_prime_1_66;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_67;
            end if;
        when square_with_reduction_special_prime_1_67 =>
            next_state <= square_with_reduction_special_prime_1_67;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_68;
            end if;
        when square_with_reduction_special_prime_1_68 =>
            next_state <= square_with_reduction_special_prime_1_68;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_69;
            end if;
        when square_with_reduction_special_prime_1_69 =>
            next_state <= square_with_reduction_special_prime_1_69;
            if(ultimate_operation = '1') then
                if(operands_size = "101") then
                    next_state <= square_with_reduction_special_prime_1_70;
                else
                    next_state <= square_with_reduction_special_prime_1_96;
                end if;
            end if;
        when square_with_reduction_special_prime_1_70 =>
            next_state <= square_with_reduction_special_prime_1_70;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_71;
            end if;
        when square_with_reduction_special_prime_1_71 =>
            next_state <= square_with_reduction_special_prime_1_71;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_72;
            end if;
        when square_with_reduction_special_prime_1_72 =>
            next_state <= square_with_reduction_special_prime_1_72;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_73;
            end if;
        when square_with_reduction_special_prime_1_73 =>
            next_state <= square_with_reduction_special_prime_1_73;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_74;
            end if;
        when square_with_reduction_special_prime_1_74 =>
            next_state <= square_with_reduction_special_prime_1_74;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_75;
            end if;
        when square_with_reduction_special_prime_1_75 =>
            next_state <= square_with_reduction_special_prime_1_75;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_76;
            end if;
        when square_with_reduction_special_prime_1_76 =>
            next_state <= square_with_reduction_special_prime_1_76;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_77;
            end if;
        when square_with_reduction_special_prime_1_77 =>
            next_state <= square_with_reduction_special_prime_1_77;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_78;
            end if;
        when square_with_reduction_special_prime_1_78 =>
            next_state <= square_with_reduction_special_prime_1_78;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_79;
            end if;
        when square_with_reduction_special_prime_1_79 =>
            next_state <= square_with_reduction_special_prime_1_79;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_80;
            end if;
        when square_with_reduction_special_prime_1_80 =>
            next_state <= square_with_reduction_special_prime_1_80;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_81;
            end if;
        when square_with_reduction_special_prime_1_81 =>
            next_state <= square_with_reduction_special_prime_1_81;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_82;
            end if;
        when square_with_reduction_special_prime_1_82 =>
            next_state <= square_with_reduction_special_prime_1_82;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_83;
            end if;
        when square_with_reduction_special_prime_1_83 =>
            next_state <= square_with_reduction_special_prime_1_83;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_84;
            end if;
        when square_with_reduction_special_prime_1_84 =>
            next_state <= square_with_reduction_special_prime_1_84;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_85;
            end if;
        when square_with_reduction_special_prime_1_85 =>
            next_state <= square_with_reduction_special_prime_1_85;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_86;
            end if;
        when square_with_reduction_special_prime_1_86 =>
            next_state <= square_with_reduction_special_prime_1_86;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_87;
            end if;
        when square_with_reduction_special_prime_1_87 =>
            next_state <= square_with_reduction_special_prime_1_87;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_88;
            end if;
        when square_with_reduction_special_prime_1_88 =>
            next_state <= square_with_reduction_special_prime_1_88;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_89;
            end if;
        when square_with_reduction_special_prime_1_89 =>
            next_state <= square_with_reduction_special_prime_1_89;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_90;
            end if;
        when square_with_reduction_special_prime_1_90 =>
            next_state <= square_with_reduction_special_prime_1_90;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_91;
            end if;
        when square_with_reduction_special_prime_1_91 =>
            next_state <= square_with_reduction_special_prime_1_91;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_92;
            end if;
        when square_with_reduction_special_prime_1_92 =>
            next_state <= square_with_reduction_special_prime_1_92;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_93;
            end if;
        when square_with_reduction_special_prime_1_93 =>
            next_state <= square_with_reduction_special_prime_1_93;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_94;
            end if;
        when square_with_reduction_special_prime_1_94 =>
            next_state <= square_with_reduction_special_prime_1_94;
            if(ultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when square_with_reduction_special_prime_1_96 =>
            next_state <= square_with_reduction_special_prime_1_96;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_97;
            end if;
        when square_with_reduction_special_prime_1_97 =>
            next_state <= square_with_reduction_special_prime_1_97;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_98;
            end if;
        when square_with_reduction_special_prime_1_98 =>
            next_state <= square_with_reduction_special_prime_1_98;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_99;
            end if;
        when square_with_reduction_special_prime_1_99 =>
            next_state <= square_with_reduction_special_prime_1_99;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_100;
            end if;
        when square_with_reduction_special_prime_1_100 =>
            next_state <= square_with_reduction_special_prime_1_100;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_101;
            end if;
        when square_with_reduction_special_prime_1_101 =>
            next_state <= square_with_reduction_special_prime_1_101;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_102;
            end if;
        when square_with_reduction_special_prime_1_102 =>
            next_state <= square_with_reduction_special_prime_1_102;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_103;
            end if;
        when square_with_reduction_special_prime_1_103 =>
            next_state <= square_with_reduction_special_prime_1_103;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_104;
            end if;
        when square_with_reduction_special_prime_1_104 =>
            next_state <= square_with_reduction_special_prime_1_104;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_105;
            end if;
        when square_with_reduction_special_prime_1_105 =>
            next_state <= square_with_reduction_special_prime_1_105;
            if(ultimate_operation = '1') then
                if(operands_size = "110") then
                    next_state <= square_with_reduction_special_prime_1_106;
                else
                    next_state <= square_with_reduction_special_prime_1_141;
                end if;
            end if;
        when square_with_reduction_special_prime_1_106 =>
            next_state <= square_with_reduction_special_prime_1_106;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_107;
            end if;
        when square_with_reduction_special_prime_1_107 =>
            next_state <= square_with_reduction_special_prime_1_107;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_108;
            end if;
        when square_with_reduction_special_prime_1_108 =>
            next_state <= square_with_reduction_special_prime_1_108;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_109;
            end if;
        when square_with_reduction_special_prime_1_109 =>
            next_state <= square_with_reduction_special_prime_1_109;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_110;
            end if;
        when square_with_reduction_special_prime_1_110 =>
            next_state <= square_with_reduction_special_prime_1_110;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_111;
            end if;
        when square_with_reduction_special_prime_1_111 =>
            next_state <= square_with_reduction_special_prime_1_111;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_112;
            end if;
        when square_with_reduction_special_prime_1_112 =>
            next_state <= square_with_reduction_special_prime_1_112;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_113;
            end if;
        when square_with_reduction_special_prime_1_113 =>
            next_state <= square_with_reduction_special_prime_1_113;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_114;
            end if;
        when square_with_reduction_special_prime_1_114 =>
            next_state <= square_with_reduction_special_prime_1_114;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_115;
            end if;
        when square_with_reduction_special_prime_1_115 =>
            next_state <= square_with_reduction_special_prime_1_115;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_116;
            end if;
        when square_with_reduction_special_prime_1_116 =>
            next_state <= square_with_reduction_special_prime_1_116;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_117;
            end if;
        when square_with_reduction_special_prime_1_117 =>
            next_state <= square_with_reduction_special_prime_1_117;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_118;
            end if;
        when square_with_reduction_special_prime_1_118 =>
            next_state <= square_with_reduction_special_prime_1_118;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_119;
            end if;
        when square_with_reduction_special_prime_1_119 =>
            next_state <= square_with_reduction_special_prime_1_119;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_120;
            end if;
        when square_with_reduction_special_prime_1_120 =>
            next_state <= square_with_reduction_special_prime_1_120;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_121;
            end if;
        when square_with_reduction_special_prime_1_121 =>
            next_state <= square_with_reduction_special_prime_1_121;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_122;
            end if;
        when square_with_reduction_special_prime_1_122 =>
            next_state <= square_with_reduction_special_prime_1_122;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_123;
            end if;
        when square_with_reduction_special_prime_1_123 =>
            next_state <= square_with_reduction_special_prime_1_123;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_124;
            end if;
        when square_with_reduction_special_prime_1_124 =>
            next_state <= square_with_reduction_special_prime_1_124;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_125;
            end if;
        when square_with_reduction_special_prime_1_125 =>
            next_state <= square_with_reduction_special_prime_1_125;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_126;
            end if;
        when square_with_reduction_special_prime_1_126 =>
            next_state <= square_with_reduction_special_prime_1_126;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_127;
            end if;
        when square_with_reduction_special_prime_1_127 =>
            next_state <= square_with_reduction_special_prime_1_127;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_128;
            end if;
        when square_with_reduction_special_prime_1_128 =>
            next_state <= square_with_reduction_special_prime_1_128;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_129;
            end if;
        when square_with_reduction_special_prime_1_129 =>
            next_state <= square_with_reduction_special_prime_1_129;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_130;
            end if;
        when square_with_reduction_special_prime_1_130 =>
            next_state <= square_with_reduction_special_prime_1_130;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_131;
            end if;
        when square_with_reduction_special_prime_1_131 =>
            next_state <= square_with_reduction_special_prime_1_131;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_132;
            end if;
        when square_with_reduction_special_prime_1_132 =>
            next_state <= square_with_reduction_special_prime_1_132;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_133;
            end if;
        when square_with_reduction_special_prime_1_133 =>
            next_state <= square_with_reduction_special_prime_1_133;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_134;
            end if;
        when square_with_reduction_special_prime_1_134 =>
            next_state <= square_with_reduction_special_prime_1_134;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_135;
            end if;
        when square_with_reduction_special_prime_1_135 =>
            next_state <= square_with_reduction_special_prime_1_135;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_136;
            end if;
        when square_with_reduction_special_prime_1_136 =>
            next_state <= square_with_reduction_special_prime_1_136;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_137;
            end if;
        when square_with_reduction_special_prime_1_137 =>
            next_state <= square_with_reduction_special_prime_1_137;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_138;
            end if;
        when square_with_reduction_special_prime_1_138 =>
            next_state <= square_with_reduction_special_prime_1_138;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_139;
            end if;
        when square_with_reduction_special_prime_1_139 =>
            next_state <= square_with_reduction_special_prime_1_139;
            if(ultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when square_with_reduction_special_prime_1_141 =>
            next_state <= square_with_reduction_special_prime_1_141;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_142;
            end if;
        when square_with_reduction_special_prime_1_142 =>
            next_state <= square_with_reduction_special_prime_1_142;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_143;
            end if;
        when square_with_reduction_special_prime_1_143 =>
            next_state <= square_with_reduction_special_prime_1_143;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_144;
            end if;
        when square_with_reduction_special_prime_1_144 =>
            next_state <= square_with_reduction_special_prime_1_144;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_145;
            end if;
        when square_with_reduction_special_prime_1_145 =>
            next_state <= square_with_reduction_special_prime_1_145;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_146;
            end if;
        when square_with_reduction_special_prime_1_146 =>
            next_state <= square_with_reduction_special_prime_1_146;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_147;
            end if;
        when square_with_reduction_special_prime_1_147 =>
            next_state <= square_with_reduction_special_prime_1_147;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_148;
            end if;
        when square_with_reduction_special_prime_1_148 =>
            next_state <= square_with_reduction_special_prime_1_148;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_149;
            end if;
        when square_with_reduction_special_prime_1_149 =>
            next_state <= square_with_reduction_special_prime_1_149;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_150;
            end if;
        when square_with_reduction_special_prime_1_150 =>
            next_state <= square_with_reduction_special_prime_1_150;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_151;
            end if;
        when square_with_reduction_special_prime_1_151 =>
            next_state <= square_with_reduction_special_prime_1_151;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_152;
            end if;
        when square_with_reduction_special_prime_1_152 =>
            next_state <= square_with_reduction_special_prime_1_152;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_153;
            end if;
        when square_with_reduction_special_prime_1_153 =>
            next_state <= square_with_reduction_special_prime_1_153;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_154;
            end if;
        when square_with_reduction_special_prime_1_154 =>
            next_state <= square_with_reduction_special_prime_1_154;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_155;
            end if;
        when square_with_reduction_special_prime_1_155 =>
            next_state <= square_with_reduction_special_prime_1_155;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_156;
            end if;
        when square_with_reduction_special_prime_1_156 =>
            next_state <= square_with_reduction_special_prime_1_156;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_157;
            end if;
        when square_with_reduction_special_prime_1_157 =>
            next_state <= square_with_reduction_special_prime_1_157;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_158;
            end if;
        when square_with_reduction_special_prime_1_158 =>
            next_state <= square_with_reduction_special_prime_1_158;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_159;
            end if;
        when square_with_reduction_special_prime_1_159 =>
            next_state <= square_with_reduction_special_prime_1_159;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_160;
            end if;
        when square_with_reduction_special_prime_1_160 =>
            next_state <= square_with_reduction_special_prime_1_160;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_161;
            end if;
        when square_with_reduction_special_prime_1_161 =>
            next_state <= square_with_reduction_special_prime_1_161;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_162;
            end if;
        when square_with_reduction_special_prime_1_162 =>
            next_state <= square_with_reduction_special_prime_1_162;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_163;
            end if;
        when square_with_reduction_special_prime_1_163 =>
            next_state <= square_with_reduction_special_prime_1_163;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_164;
            end if;
        when square_with_reduction_special_prime_1_164 =>
            next_state <= square_with_reduction_special_prime_1_164;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_165;
            end if;
        when square_with_reduction_special_prime_1_165 =>
            next_state <= square_with_reduction_special_prime_1_165;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_166;
            end if;
        when square_with_reduction_special_prime_1_166 =>
            next_state <= square_with_reduction_special_prime_1_166;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_167;
            end if;
        when square_with_reduction_special_prime_1_167 =>
            next_state <= square_with_reduction_special_prime_1_167;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_168;
            end if;
        when square_with_reduction_special_prime_1_168 =>
            next_state <= square_with_reduction_special_prime_1_168;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_169;
            end if;
        when square_with_reduction_special_prime_1_169 =>
            next_state <= square_with_reduction_special_prime_1_169;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_170;
            end if;
        when square_with_reduction_special_prime_1_170 =>
            next_state <= square_with_reduction_special_prime_1_170;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_171;
            end if;
        when square_with_reduction_special_prime_1_171 =>
            next_state <= square_with_reduction_special_prime_1_171;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_172;
            end if;
        when square_with_reduction_special_prime_1_172 =>
            next_state <= square_with_reduction_special_prime_1_172;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_173;
            end if;
        when square_with_reduction_special_prime_1_173 =>
            next_state <= square_with_reduction_special_prime_1_173;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_174;
            end if;
        when square_with_reduction_special_prime_1_174 =>
            next_state <= square_with_reduction_special_prime_1_174;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_175;
            end if;
        when square_with_reduction_special_prime_1_175 =>
            next_state <= square_with_reduction_special_prime_1_175;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_176;
            end if;
        when square_with_reduction_special_prime_1_176 =>
            next_state <= square_with_reduction_special_prime_1_176;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_177;
            end if;
        when square_with_reduction_special_prime_1_177 =>
            next_state <= square_with_reduction_special_prime_1_177;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_178;
            end if;
        when square_with_reduction_special_prime_1_178 =>
            next_state <= square_with_reduction_special_prime_1_178;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_179;
            end if;
        when square_with_reduction_special_prime_1_179 =>
            next_state <= square_with_reduction_special_prime_1_179;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_180;
            end if;
        when square_with_reduction_special_prime_1_180 =>
            next_state <= square_with_reduction_special_prime_1_180;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_181;
            end if;
        when square_with_reduction_special_prime_1_181 =>
            next_state <= square_with_reduction_special_prime_1_181;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_182;
            end if;
        when square_with_reduction_special_prime_1_182 =>
            next_state <= square_with_reduction_special_prime_1_182;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_183;
            end if;
        when square_with_reduction_special_prime_1_183 =>
            next_state <= square_with_reduction_special_prime_1_183;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_184;
            end if;
        when square_with_reduction_special_prime_1_184 =>
            next_state <= square_with_reduction_special_prime_1_184;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_185;
            end if;
        when square_with_reduction_special_prime_1_185 =>
            next_state <= square_with_reduction_special_prime_1_185;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_186;
            end if;
        when square_with_reduction_special_prime_1_186 =>
            next_state <= square_with_reduction_special_prime_1_186;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_187;
            end if;
        when square_with_reduction_special_prime_1_187 =>
            next_state <= square_with_reduction_special_prime_1_187;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_188;
            end if;
        when square_with_reduction_special_prime_1_188 =>
            next_state <= square_with_reduction_special_prime_1_188;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_189;
            end if;
        when square_with_reduction_special_prime_1_189 =>
            next_state <= square_with_reduction_special_prime_1_189;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_190;
            end if;
        when square_with_reduction_special_prime_1_190 =>
            next_state <= square_with_reduction_special_prime_1_190;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_191;
            end if;
        when square_with_reduction_special_prime_1_191 =>
            next_state <= square_with_reduction_special_prime_1_191;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_192;
            end if;
        when square_with_reduction_special_prime_1_192 =>
            next_state <= square_with_reduction_special_prime_1_192;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_193;
            end if;
        when square_with_reduction_special_prime_1_193 =>
            next_state <= square_with_reduction_special_prime_1_193;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_194;
            end if;
        when square_with_reduction_special_prime_1_194 =>
            next_state <= square_with_reduction_special_prime_1_194;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_195;
            end if;
        when square_with_reduction_special_prime_1_195 =>
            next_state <= square_with_reduction_special_prime_1_195;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1_196;
            end if;
        when square_with_reduction_special_prime_1_196 =>
            next_state <= square_with_reduction_special_prime_1_196;
            if(ultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when square_with_reduction_special_prime_2_0 => 
            next_state <= square_with_reduction_special_prime_2_0;
            if(ultimate_operation = '1') then
                if(operands_size = "001") then
                    next_state <= square_with_reduction_special_prime_2_1;
                else
                    next_state <= square_with_reduction_special_prime_2_4;
                end if;
            end if;
            
        when square_with_reduction_special_prime_2_1 => 
            next_state <= square_with_reduction_special_prime_2_1;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_2;
            end if;
        when square_with_reduction_special_prime_2_2 => 
            next_state <= square_with_reduction_special_prime_2_2;
            if(ultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when square_with_reduction_special_prime_2_4 => 
            next_state <= square_with_reduction_special_prime_2_4;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_5;
            end if;
        when square_with_reduction_special_prime_2_5 => 
            next_state <= square_with_reduction_special_prime_2_5;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_6;
            end if;
        when square_with_reduction_special_prime_2_6 => 
            next_state <= square_with_reduction_special_prime_2_6;
            if(ultimate_operation = '1') then
                if(operands_size = "010") then
                    next_state <= square_with_reduction_special_prime_2_7;
                else
                    next_state <= square_with_reduction_special_prime_2_13;
                end if;
            end if;
        when square_with_reduction_special_prime_2_7 =>
            next_state <= square_with_reduction_special_prime_2_7;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_8;
            end if;
        when square_with_reduction_special_prime_2_8 =>
            next_state <= square_with_reduction_special_prime_2_8;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_9;
            end if;
        when square_with_reduction_special_prime_2_9 =>
            next_state <= square_with_reduction_special_prime_2_9;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_10;
            end if;
        when square_with_reduction_special_prime_2_10 =>
            next_state <= square_with_reduction_special_prime_2_10;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_11;
            end if;
        when square_with_reduction_special_prime_2_11 =>
            next_state <= square_with_reduction_special_prime_2_11;
            if(ultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when square_with_reduction_special_prime_2_13 => 
            next_state <= square_with_reduction_special_prime_2_13;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_14;
            end if;
        when square_with_reduction_special_prime_2_14 => 
            next_state <= square_with_reduction_special_prime_2_14;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_15;
            end if;
        when square_with_reduction_special_prime_2_15 => 
            next_state <= square_with_reduction_special_prime_2_15;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_16;
            end if;
        when square_with_reduction_special_prime_2_16 => 
            next_state <= square_with_reduction_special_prime_2_16;
            if(ultimate_operation = '1') then
                if(operands_size = "011") then
                    next_state <= square_with_reduction_special_prime_2_17;
                else
                    next_state <= square_with_reduction_special_prime_2_28;
                end if;
            end if;
        when square_with_reduction_special_prime_2_17 =>
            next_state <= square_with_reduction_special_prime_2_17;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_18;
            end if;
        when square_with_reduction_special_prime_2_18 =>
            next_state <= square_with_reduction_special_prime_2_18;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_19;
            end if;
        when square_with_reduction_special_prime_2_19 =>
            next_state <= square_with_reduction_special_prime_2_19;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_20;
            end if;
        when square_with_reduction_special_prime_2_20 =>
            next_state <= square_with_reduction_special_prime_2_20;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_21;
            end if;
        when square_with_reduction_special_prime_2_21 =>
            next_state <= square_with_reduction_special_prime_2_21;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_22;
            end if;
        when square_with_reduction_special_prime_2_22 =>
            next_state <= square_with_reduction_special_prime_2_22;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_23;
            end if;
        when square_with_reduction_special_prime_2_23 =>
            next_state <= square_with_reduction_special_prime_2_23;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_24;
            end if;
        when square_with_reduction_special_prime_2_24 =>
            next_state <= square_with_reduction_special_prime_2_24;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_25;
            end if;
        when square_with_reduction_special_prime_2_25 =>
            next_state <= square_with_reduction_special_prime_2_25;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_26;
            end if;
        when square_with_reduction_special_prime_2_26 =>
            next_state <= square_with_reduction_special_prime_2_26;
            if(ultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when square_with_reduction_special_prime_2_28 => 
            next_state <= square_with_reduction_special_prime_2_28;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_29;
            end if;
        when square_with_reduction_special_prime_2_29 => 
            next_state <= square_with_reduction_special_prime_2_29;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_30;
            end if;
        when square_with_reduction_special_prime_2_30 => 
            next_state <= square_with_reduction_special_prime_2_30;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_31;
            end if;
        when square_with_reduction_special_prime_2_31 => 
            next_state <= square_with_reduction_special_prime_2_31;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_32;
            end if;
        when square_with_reduction_special_prime_2_32 => 
            next_state <= square_with_reduction_special_prime_2_32;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_33;
            end if;
        when square_with_reduction_special_prime_2_33 => 
            next_state <= square_with_reduction_special_prime_2_33;
            if(ultimate_operation = '1') then
                if(operands_size = "100") then
                    next_state <= square_with_reduction_special_prime_2_34;
                else
                    next_state <= square_with_reduction_special_prime_2_51;
                end if;
            end if;
        when square_with_reduction_special_prime_2_34 => 
            next_state <= square_with_reduction_special_prime_2_34;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_35;
            end if;
        when square_with_reduction_special_prime_2_35 => 
            next_state <= square_with_reduction_special_prime_2_35;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_36;
            end if;
        when square_with_reduction_special_prime_2_36 => 
            next_state <= square_with_reduction_special_prime_2_36;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_37;
            end if;
        when square_with_reduction_special_prime_2_37 => 
            next_state <= square_with_reduction_special_prime_2_37;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_38;
            end if;
        when square_with_reduction_special_prime_2_38 => 
            next_state <= square_with_reduction_special_prime_2_38;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_39;
            end if;
        when square_with_reduction_special_prime_2_39 => 
            next_state <= square_with_reduction_special_prime_2_39;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_40;
            end if;
        when square_with_reduction_special_prime_2_40 => 
            next_state <= square_with_reduction_special_prime_2_40;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_41;
            end if;
        when square_with_reduction_special_prime_2_41 => 
            next_state <= square_with_reduction_special_prime_2_41;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_42;
            end if;
        when square_with_reduction_special_prime_2_42 => 
            next_state <= square_with_reduction_special_prime_2_42;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_43;
            end if;
        when square_with_reduction_special_prime_2_43 => 
            next_state <= square_with_reduction_special_prime_2_43;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_44;
            end if;
        when square_with_reduction_special_prime_2_44 => 
            next_state <= square_with_reduction_special_prime_2_44;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_45;
            end if;
        when square_with_reduction_special_prime_2_45 => 
            next_state <= square_with_reduction_special_prime_2_45;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_46;
            end if;
        when square_with_reduction_special_prime_2_46 => 
            next_state <= square_with_reduction_special_prime_2_46;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_47;
            end if;
        when square_with_reduction_special_prime_2_47 => 
            next_state <= square_with_reduction_special_prime_2_47;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_48;
            end if;
        when square_with_reduction_special_prime_2_48 => 
            next_state <= square_with_reduction_special_prime_2_48;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_49;
            end if;
        when square_with_reduction_special_prime_2_49 => 
            next_state <= square_with_reduction_special_prime_2_49;
            if(ultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when square_with_reduction_special_prime_2_51 => 
            next_state <= square_with_reduction_special_prime_2_51;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_52;
            end if;
        when square_with_reduction_special_prime_2_52 => 
            next_state <= square_with_reduction_special_prime_2_52;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_53;
            end if;
        when square_with_reduction_special_prime_2_53 => 
            next_state <= square_with_reduction_special_prime_2_53;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_54;
            end if;
        when square_with_reduction_special_prime_2_54 => 
            next_state <= square_with_reduction_special_prime_2_54;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_55;
            end if;
        when square_with_reduction_special_prime_2_55 => 
            next_state <= square_with_reduction_special_prime_2_55;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_56;
            end if;
        when square_with_reduction_special_prime_2_56 => 
            next_state <= square_with_reduction_special_prime_2_56;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_57;
            end if;
        when square_with_reduction_special_prime_2_57 => 
            next_state <= square_with_reduction_special_prime_2_57;
            if(ultimate_operation = '1') then
                if(operands_size = "101") then
                    next_state <= square_with_reduction_special_prime_2_58;
                else
                    next_state <= square_with_reduction_special_prime_2_83;
                end if;
            end if;
        when square_with_reduction_special_prime_2_58 => 
            next_state <= square_with_reduction_special_prime_2_58;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_59;
            end if;
        when square_with_reduction_special_prime_2_59 => 
            next_state <= square_with_reduction_special_prime_2_59;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_60;
            end if;
        when square_with_reduction_special_prime_2_60 => 
            next_state <= square_with_reduction_special_prime_2_60;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_61;
            end if;
        when square_with_reduction_special_prime_2_61 => 
            next_state <= square_with_reduction_special_prime_2_61;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_62;
            end if;
        when square_with_reduction_special_prime_2_62 => 
            next_state <= square_with_reduction_special_prime_2_62;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_63;
            end if;
        when square_with_reduction_special_prime_2_63 => 
            next_state <= square_with_reduction_special_prime_2_63;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_64;
            end if;
        when square_with_reduction_special_prime_2_64 => 
            next_state <= square_with_reduction_special_prime_2_64;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_65;
            end if;
        when square_with_reduction_special_prime_2_65 => 
            next_state <= square_with_reduction_special_prime_2_65;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_66;
            end if;
        when square_with_reduction_special_prime_2_66 => 
            next_state <= square_with_reduction_special_prime_2_66;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_67;
            end if;
        when square_with_reduction_special_prime_2_67 => 
            next_state <= square_with_reduction_special_prime_2_67;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_68;
            end if;
        when square_with_reduction_special_prime_2_68 => 
            next_state <= square_with_reduction_special_prime_2_68;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_69;
            end if;
        when square_with_reduction_special_prime_2_69 => 
            next_state <= square_with_reduction_special_prime_2_69;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_70;
            end if;
        when square_with_reduction_special_prime_2_70 => 
            next_state <= square_with_reduction_special_prime_2_70;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_71;
            end if;
        when square_with_reduction_special_prime_2_71 => 
            next_state <= square_with_reduction_special_prime_2_71;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_72;
            end if;
        when square_with_reduction_special_prime_2_72 => 
            next_state <= square_with_reduction_special_prime_2_72;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_73;
            end if;
        when square_with_reduction_special_prime_2_73 => 
            next_state <= square_with_reduction_special_prime_2_73;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_74;
            end if;
        when square_with_reduction_special_prime_2_74 => 
            next_state <= square_with_reduction_special_prime_2_74;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_75;
            end if;
        when square_with_reduction_special_prime_2_75 => 
            next_state <= square_with_reduction_special_prime_2_75;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_76;
            end if;
        when square_with_reduction_special_prime_2_76 => 
            next_state <= square_with_reduction_special_prime_2_76;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_77;
            end if;
        when square_with_reduction_special_prime_2_77 => 
            next_state <= square_with_reduction_special_prime_2_77;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_78;
            end if;
        when square_with_reduction_special_prime_2_78 => 
            next_state <= square_with_reduction_special_prime_2_78;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_79;
            end if;
        when square_with_reduction_special_prime_2_79 => 
            next_state <= square_with_reduction_special_prime_2_79;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_80;
            end if;
        when square_with_reduction_special_prime_2_80 => 
            next_state <= square_with_reduction_special_prime_2_80;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_81;
            end if;
        when square_with_reduction_special_prime_2_81 => 
            next_state <= square_with_reduction_special_prime_2_81;
            if(ultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when square_with_reduction_special_prime_2_83 =>
            next_state <= square_with_reduction_special_prime_2_83;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_84;
            end if;
        when square_with_reduction_special_prime_2_84 =>
            next_state <= square_with_reduction_special_prime_2_84;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_85;
            end if;
        when square_with_reduction_special_prime_2_85 =>
            next_state <= square_with_reduction_special_prime_2_85;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_86;
            end if;
        when square_with_reduction_special_prime_2_86 =>
            next_state <= square_with_reduction_special_prime_2_86;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_87;
            end if;
        when square_with_reduction_special_prime_2_87 =>
            next_state <= square_with_reduction_special_prime_2_87;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_88;
            end if;
        when square_with_reduction_special_prime_2_88 =>
            next_state <= square_with_reduction_special_prime_2_88;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_89;
            end if;
        when square_with_reduction_special_prime_2_89 =>
            next_state <= square_with_reduction_special_prime_2_89;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_90;
            end if;
        when square_with_reduction_special_prime_2_90 =>
            next_state <= square_with_reduction_special_prime_2_90;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_91;
            end if;
        when square_with_reduction_special_prime_2_91 =>
            next_state <= square_with_reduction_special_prime_2_91;
            if(ultimate_operation = '1') then
                if(operands_size = "110") then
                    next_state <= square_with_reduction_special_prime_2_92;
                else
                    next_state <= square_with_reduction_special_prime_2_126;
                end if;
            end if;
        when square_with_reduction_special_prime_2_92 =>
            next_state <= square_with_reduction_special_prime_2_92;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_93;
            end if;
        when square_with_reduction_special_prime_2_93 =>
            next_state <= square_with_reduction_special_prime_2_93;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_94;
            end if;
        when square_with_reduction_special_prime_2_94 =>
            next_state <= square_with_reduction_special_prime_2_94;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_95;
            end if;
        when square_with_reduction_special_prime_2_95 =>
            next_state <= square_with_reduction_special_prime_2_95;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_96;
            end if;
        when square_with_reduction_special_prime_2_96 =>
            next_state <= square_with_reduction_special_prime_2_96;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_97;
            end if;
        when square_with_reduction_special_prime_2_97 =>
            next_state <= square_with_reduction_special_prime_2_97;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_98;
            end if;
        when square_with_reduction_special_prime_2_98 =>
            next_state <= square_with_reduction_special_prime_2_98;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_99;
            end if;
        when square_with_reduction_special_prime_2_99 =>
            next_state <= square_with_reduction_special_prime_2_99;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_100;
            end if;
        when square_with_reduction_special_prime_2_100 =>
            next_state <= square_with_reduction_special_prime_2_100;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_101;
            end if;
        when square_with_reduction_special_prime_2_101 =>
            next_state <= square_with_reduction_special_prime_2_101;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_102;
            end if;
        when square_with_reduction_special_prime_2_102 =>
            next_state <= square_with_reduction_special_prime_2_102;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_103;
            end if;
        when square_with_reduction_special_prime_2_103 =>
            next_state <= square_with_reduction_special_prime_2_103;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_104;
            end if;
        when square_with_reduction_special_prime_2_104 =>
            next_state <= square_with_reduction_special_prime_2_104;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_105;
            end if;
        when square_with_reduction_special_prime_2_105 =>
            next_state <= square_with_reduction_special_prime_2_105;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_106;
            end if;
        when square_with_reduction_special_prime_2_106 =>
            next_state <= square_with_reduction_special_prime_2_106;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_107;
            end if;
        when square_with_reduction_special_prime_2_107 =>
            next_state <= square_with_reduction_special_prime_2_107;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_108;
            end if;
        when square_with_reduction_special_prime_2_108 =>
            next_state <= square_with_reduction_special_prime_2_108;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_109;
            end if;
        when square_with_reduction_special_prime_2_109 =>
            next_state <= square_with_reduction_special_prime_2_109;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_110;
            end if;
        when square_with_reduction_special_prime_2_110 =>
            next_state <= square_with_reduction_special_prime_2_110;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_111;
            end if;
        when square_with_reduction_special_prime_2_111 =>
            next_state <= square_with_reduction_special_prime_2_111;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_112;
            end if;
        when square_with_reduction_special_prime_2_112 =>
            next_state <= square_with_reduction_special_prime_2_112;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_113;
            end if;
        when square_with_reduction_special_prime_2_113 =>
            next_state <= square_with_reduction_special_prime_2_113;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_114;
            end if;
        when square_with_reduction_special_prime_2_114 =>
            next_state <= square_with_reduction_special_prime_2_114;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_115;
            end if;
        when square_with_reduction_special_prime_2_115 =>
            next_state <= square_with_reduction_special_prime_2_115;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_116;
            end if;
        when square_with_reduction_special_prime_2_116 =>
            next_state <= square_with_reduction_special_prime_2_116;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_117;
            end if;
        when square_with_reduction_special_prime_2_117 =>
            next_state <= square_with_reduction_special_prime_2_117;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_118;
            end if;
        when square_with_reduction_special_prime_2_118 =>
            next_state <= square_with_reduction_special_prime_2_118;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_119;
            end if;
        when square_with_reduction_special_prime_2_119 =>
            next_state <= square_with_reduction_special_prime_2_119;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_120;
            end if;
        when square_with_reduction_special_prime_2_120 =>
            next_state <= square_with_reduction_special_prime_2_120;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_121;
            end if;
        when square_with_reduction_special_prime_2_121 =>
            next_state <= square_with_reduction_special_prime_2_121;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_122;
            end if;
        when square_with_reduction_special_prime_2_122 =>
            next_state <= square_with_reduction_special_prime_2_122;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_123;
            end if;
        when square_with_reduction_special_prime_2_123 =>
            next_state <= square_with_reduction_special_prime_2_123;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_124;
            end if;
        when square_with_reduction_special_prime_2_124 =>
            next_state <= square_with_reduction_special_prime_2_124;
            if(ultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when square_with_reduction_special_prime_2_126 =>
            next_state <= square_with_reduction_special_prime_2_126;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_127;
            end if;
        when square_with_reduction_special_prime_2_127 =>
            next_state <= square_with_reduction_special_prime_2_127;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_128;
            end if;
        when square_with_reduction_special_prime_2_128 =>
            next_state <= square_with_reduction_special_prime_2_128;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_129;
            end if;
        when square_with_reduction_special_prime_2_129 =>
            next_state <= square_with_reduction_special_prime_2_129;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_130;
            end if;
        when square_with_reduction_special_prime_2_130 =>
            next_state <= square_with_reduction_special_prime_2_130;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_131;
            end if;
        when square_with_reduction_special_prime_2_131 =>
            next_state <= square_with_reduction_special_prime_2_131;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_132;
            end if;
        when square_with_reduction_special_prime_2_132 =>
            next_state <= square_with_reduction_special_prime_2_132;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_133;
            end if;
        when square_with_reduction_special_prime_2_133 =>
            next_state <= square_with_reduction_special_prime_2_133;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_134;
            end if;
        when square_with_reduction_special_prime_2_134 =>
            next_state <= square_with_reduction_special_prime_2_134;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_135;
            end if;
        when square_with_reduction_special_prime_2_135 =>
            next_state <= square_with_reduction_special_prime_2_135;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_136;
            end if;
        when square_with_reduction_special_prime_2_136 =>
            next_state <= square_with_reduction_special_prime_2_136;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_137;
            end if;
        when square_with_reduction_special_prime_2_137 =>
            next_state <= square_with_reduction_special_prime_2_137;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_138;
            end if;
        when square_with_reduction_special_prime_2_138 =>
            next_state <= square_with_reduction_special_prime_2_138;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_139;
            end if;
        when square_with_reduction_special_prime_2_139 =>
            next_state <= square_with_reduction_special_prime_2_139;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_140;
            end if;
        when square_with_reduction_special_prime_2_140 =>
            next_state <= square_with_reduction_special_prime_2_140;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_141;
            end if;
        when square_with_reduction_special_prime_2_141 =>
            next_state <= square_with_reduction_special_prime_2_141;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_142;
            end if;
        when square_with_reduction_special_prime_2_142 =>
            next_state <= square_with_reduction_special_prime_2_142;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_143;
            end if;
        when square_with_reduction_special_prime_2_143 =>
            next_state <= square_with_reduction_special_prime_2_143;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_144;
            end if;
        when square_with_reduction_special_prime_2_144 =>
            next_state <= square_with_reduction_special_prime_2_144;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_145;
            end if;
        when square_with_reduction_special_prime_2_145 =>
            next_state <= square_with_reduction_special_prime_2_145;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_146;
            end if;
        when square_with_reduction_special_prime_2_146 =>
            next_state <= square_with_reduction_special_prime_2_146;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_147;
            end if;
        when square_with_reduction_special_prime_2_147 =>
            next_state <= square_with_reduction_special_prime_2_147;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_148;
            end if;
        when square_with_reduction_special_prime_2_148 =>
            next_state <= square_with_reduction_special_prime_2_148;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_149;
            end if;
        when square_with_reduction_special_prime_2_149 =>
            next_state <= square_with_reduction_special_prime_2_149;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_150;
            end if;
        when square_with_reduction_special_prime_2_150 =>
            next_state <= square_with_reduction_special_prime_2_150;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_151;
            end if;
        when square_with_reduction_special_prime_2_151 =>
            next_state <= square_with_reduction_special_prime_2_151;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_152;
            end if;
        when square_with_reduction_special_prime_2_152 =>
            next_state <= square_with_reduction_special_prime_2_152;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_153;
            end if;
        when square_with_reduction_special_prime_2_153 =>
            next_state <= square_with_reduction_special_prime_2_153;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_154;
            end if;
        when square_with_reduction_special_prime_2_154 =>
            next_state <= square_with_reduction_special_prime_2_154;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_155;
            end if;
        when square_with_reduction_special_prime_2_155 =>
            next_state <= square_with_reduction_special_prime_2_155;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_156;
            end if;
        when square_with_reduction_special_prime_2_156 =>
            next_state <= square_with_reduction_special_prime_2_156;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_157;
            end if;
        when square_with_reduction_special_prime_2_157 =>
            next_state <= square_with_reduction_special_prime_2_157;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_158;
            end if;
        when square_with_reduction_special_prime_2_158 =>
            next_state <= square_with_reduction_special_prime_2_158;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_159;
            end if;
        when square_with_reduction_special_prime_2_159 =>
            next_state <= square_with_reduction_special_prime_2_159;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_160;
            end if;
        when square_with_reduction_special_prime_2_160 =>
            next_state <= square_with_reduction_special_prime_2_160;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_161;
            end if;
        when square_with_reduction_special_prime_2_161 =>
            next_state <= square_with_reduction_special_prime_2_161;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_162;
            end if;
        when square_with_reduction_special_prime_2_162 =>
            next_state <= square_with_reduction_special_prime_2_162;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_163;
            end if;
        when square_with_reduction_special_prime_2_163 =>
            next_state <= square_with_reduction_special_prime_2_163;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_164;
            end if;
        when square_with_reduction_special_prime_2_164 =>
            next_state <= square_with_reduction_special_prime_2_164;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_165;
            end if;
        when square_with_reduction_special_prime_2_165 =>
            next_state <= square_with_reduction_special_prime_2_165;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_166;
            end if;
        when square_with_reduction_special_prime_2_166 =>
            next_state <= square_with_reduction_special_prime_2_166;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_167;
            end if;
        when square_with_reduction_special_prime_2_167 =>
            next_state <= square_with_reduction_special_prime_2_167;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_168;
            end if;
        when square_with_reduction_special_prime_2_168 =>
            next_state <= square_with_reduction_special_prime_2_168;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_169;
            end if;
        when square_with_reduction_special_prime_2_169 =>
            next_state <= square_with_reduction_special_prime_2_169;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_170;
            end if;
        when square_with_reduction_special_prime_2_170 =>
            next_state <= square_with_reduction_special_prime_2_170;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_171;
            end if;
        when square_with_reduction_special_prime_2_171 =>
            next_state <= square_with_reduction_special_prime_2_171;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_172;
            end if;
        when square_with_reduction_special_prime_2_172 =>
            next_state <= square_with_reduction_special_prime_2_172;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_173;
            end if;
        when square_with_reduction_special_prime_2_173 =>
            next_state <= square_with_reduction_special_prime_2_173;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_174;
            end if;
        when square_with_reduction_special_prime_2_174 =>
            next_state <= square_with_reduction_special_prime_2_174;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_175;
            end if;
        when square_with_reduction_special_prime_2_175 =>
            next_state <= square_with_reduction_special_prime_2_175;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_176;
            end if;
        when square_with_reduction_special_prime_2_176 =>
            next_state <= square_with_reduction_special_prime_2_176;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_177;
            end if;
        when square_with_reduction_special_prime_2_177 =>
            next_state <= square_with_reduction_special_prime_2_177;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_178;
            end if;
        when square_with_reduction_special_prime_2_178 =>
            next_state <= square_with_reduction_special_prime_2_178;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_2_179;
            end if;
        when square_with_reduction_special_prime_2_179 =>
            next_state <= square_with_reduction_special_prime_2_179;
            if(ultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when square_with_reduction_special_prime_3_0 => 
            next_state <= square_with_reduction_special_prime_3_0;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_1;
            end if;
        when square_with_reduction_special_prime_3_1 => 
            next_state <= square_with_reduction_special_prime_3_1;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_2;
            end if;
        when square_with_reduction_special_prime_3_2 => 
            next_state <= square_with_reduction_special_prime_3_2;
            if(ultimate_operation = '1') then
                if(operands_size = "010") then
                    next_state <= square_with_reduction_special_prime_3_3;
                else
                    next_state <= square_with_reduction_special_prime_3_7;
                end if;
            end if;
        when square_with_reduction_special_prime_3_3 =>
            next_state <= square_with_reduction_special_prime_3_3;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_4;
            end if;
        when square_with_reduction_special_prime_3_4 =>
            next_state <= square_with_reduction_special_prime_3_4;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_5;
            end if;
        when square_with_reduction_special_prime_3_5 =>
            next_state <= square_with_reduction_special_prime_3_5;
            if(ultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when square_with_reduction_special_prime_3_7 => 
            next_state <= square_with_reduction_special_prime_3_7;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_8;
            end if;
        when square_with_reduction_special_prime_3_8 => 
            next_state <= square_with_reduction_special_prime_3_8;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_9;
            end if;
        when square_with_reduction_special_prime_3_9 => 
            next_state <= square_with_reduction_special_prime_3_9;
            if(ultimate_operation = '1') then
                if(operands_size = "011") then
                    next_state <= square_with_reduction_special_prime_3_10;
                else
                    next_state <= square_with_reduction_special_prime_3_19;
                end if;
            end if;
        when square_with_reduction_special_prime_3_10 =>
            next_state <= square_with_reduction_special_prime_3_10;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_11;
            end if;
        when square_with_reduction_special_prime_3_11 =>
            next_state <= square_with_reduction_special_prime_3_11;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_12;
            end if;
        when square_with_reduction_special_prime_3_12 =>
            next_state <= square_with_reduction_special_prime_3_12;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_13;
            end if;
        when square_with_reduction_special_prime_3_13 =>
            next_state <= square_with_reduction_special_prime_3_13;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_14;
            end if;
        when square_with_reduction_special_prime_3_14 =>
            next_state <= square_with_reduction_special_prime_3_14;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_15;
            end if;
        when square_with_reduction_special_prime_3_15 =>
            next_state <= square_with_reduction_special_prime_3_15;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_16;
            end if;
        when square_with_reduction_special_prime_3_16 =>
            next_state <= square_with_reduction_special_prime_3_16;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_17;
            end if;
        when square_with_reduction_special_prime_3_17 =>
            next_state <= square_with_reduction_special_prime_3_17;
            if(ultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when square_with_reduction_special_prime_3_19 => 
            next_state <= square_with_reduction_special_prime_3_19;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_20;
            end if;
        when square_with_reduction_special_prime_3_20 => 
            next_state <= square_with_reduction_special_prime_3_20;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_21;
            end if;
        when square_with_reduction_special_prime_3_21 => 
            next_state <= square_with_reduction_special_prime_3_21;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_22;
            end if;
        when square_with_reduction_special_prime_3_22 => 
            next_state <= square_with_reduction_special_prime_3_22;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_23;
            end if;
        when square_with_reduction_special_prime_3_23 => 
            next_state <= square_with_reduction_special_prime_3_23;
            if(ultimate_operation = '1') then
                if(operands_size = "100") then
                    next_state <= square_with_reduction_special_prime_3_24;
                else
                    next_state <= square_with_reduction_special_prime_3_39;
                end if;
            end if;
        when square_with_reduction_special_prime_3_24 =>
            next_state <= square_with_reduction_special_prime_3_24;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_25;
            end if;
        when square_with_reduction_special_prime_3_25 =>
            next_state <= square_with_reduction_special_prime_3_25;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_26;
            end if;
        when square_with_reduction_special_prime_3_26 =>
            next_state <= square_with_reduction_special_prime_3_26;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_27;
            end if;
        when square_with_reduction_special_prime_3_27 =>
            next_state <= square_with_reduction_special_prime_3_27;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_28;
            end if;
        when square_with_reduction_special_prime_3_28 =>
            next_state <= square_with_reduction_special_prime_3_28;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_29;
            end if;
        when square_with_reduction_special_prime_3_29 =>
            next_state <= square_with_reduction_special_prime_3_29;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_30;
            end if;
        when square_with_reduction_special_prime_3_30 =>
            next_state <= square_with_reduction_special_prime_3_30;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_31;
            end if;
        when square_with_reduction_special_prime_3_31 =>
            next_state <= square_with_reduction_special_prime_3_31;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_32;
            end if;
        when square_with_reduction_special_prime_3_32 =>
            next_state <= square_with_reduction_special_prime_3_32;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_33;
            end if;
        when square_with_reduction_special_prime_3_33 =>
            next_state <= square_with_reduction_special_prime_3_33;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_34;
            end if;
        when square_with_reduction_special_prime_3_34 =>
            next_state <= square_with_reduction_special_prime_3_34;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_35;
            end if;
        when square_with_reduction_special_prime_3_35 =>
            next_state <= square_with_reduction_special_prime_3_35;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_36;
            end if;
        when square_with_reduction_special_prime_3_36 =>
            next_state <= square_with_reduction_special_prime_3_36;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_37;
            end if;
        when square_with_reduction_special_prime_3_37 =>
            next_state <= square_with_reduction_special_prime_3_37;
            if(ultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when square_with_reduction_special_prime_3_39 => 
            next_state <= square_with_reduction_special_prime_3_39;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_40;
            end if;
        when square_with_reduction_special_prime_3_40 => 
            next_state <= square_with_reduction_special_prime_3_40;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_41;
            end if;
        when square_with_reduction_special_prime_3_41 => 
            next_state <= square_with_reduction_special_prime_3_41;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_42;
            end if;
        when square_with_reduction_special_prime_3_42 => 
            next_state <= square_with_reduction_special_prime_3_42;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_43;
            end if;
        when square_with_reduction_special_prime_3_43 => 
            next_state <= square_with_reduction_special_prime_3_43;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_44;
            end if;
        when square_with_reduction_special_prime_3_44 => 
            next_state <= square_with_reduction_special_prime_3_44;
            if(ultimate_operation = '1') then
                if(operands_size = "101") then
                    next_state <= square_with_reduction_special_prime_3_45;
                else
                    next_state <= square_with_reduction_special_prime_3_68;
                end if;
            end if;
        when square_with_reduction_special_prime_3_45 =>
            next_state <= square_with_reduction_special_prime_3_45;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_46;
            end if;
        when square_with_reduction_special_prime_3_46 =>
            next_state <= square_with_reduction_special_prime_3_46;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_47;
            end if;
        when square_with_reduction_special_prime_3_47 =>
            next_state <= square_with_reduction_special_prime_3_47;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_48;
            end if;
        when square_with_reduction_special_prime_3_48 =>
            next_state <= square_with_reduction_special_prime_3_48;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_49;
            end if;
        when square_with_reduction_special_prime_3_49 =>
            next_state <= square_with_reduction_special_prime_3_49;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_50;
            end if;
        when square_with_reduction_special_prime_3_50 =>
            next_state <= square_with_reduction_special_prime_3_50;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_51;
            end if;
        when square_with_reduction_special_prime_3_51 =>
            next_state <= square_with_reduction_special_prime_3_51;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_52;
            end if;
        when square_with_reduction_special_prime_3_52 =>
            next_state <= square_with_reduction_special_prime_3_52;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_53;
            end if;
        when square_with_reduction_special_prime_3_53 =>
            next_state <= square_with_reduction_special_prime_3_53;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_54;
            end if;
        when square_with_reduction_special_prime_3_54 =>
            next_state <= square_with_reduction_special_prime_3_54;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_55;
            end if;
        when square_with_reduction_special_prime_3_55 =>
            next_state <= square_with_reduction_special_prime_3_55;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_56;
            end if;
        when square_with_reduction_special_prime_3_56 =>
            next_state <= square_with_reduction_special_prime_3_56;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_57;
            end if;
        when square_with_reduction_special_prime_3_57 =>
            next_state <= square_with_reduction_special_prime_3_57;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_58;
            end if;
        when square_with_reduction_special_prime_3_58 =>
            next_state <= square_with_reduction_special_prime_3_58;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_59;
            end if;
        when square_with_reduction_special_prime_3_59 =>
            next_state <= square_with_reduction_special_prime_3_59;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_60;
            end if;
        when square_with_reduction_special_prime_3_60 =>
            next_state <= square_with_reduction_special_prime_3_60;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_61;
            end if;
        when square_with_reduction_special_prime_3_61 =>
            next_state <= square_with_reduction_special_prime_3_61;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_62;
            end if;
        when square_with_reduction_special_prime_3_62 =>
            next_state <= square_with_reduction_special_prime_3_62;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_63;
            end if;
        when square_with_reduction_special_prime_3_63 =>
            next_state <= square_with_reduction_special_prime_3_63;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_64;
            end if;
        when square_with_reduction_special_prime_3_64 =>
            next_state <= square_with_reduction_special_prime_3_64;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_65;
            end if;
        when square_with_reduction_special_prime_3_65 =>
            next_state <= square_with_reduction_special_prime_3_65;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_66;
            end if;
        when square_with_reduction_special_prime_3_66 =>
            next_state <= square_with_reduction_special_prime_3_66;
            if(ultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when square_with_reduction_special_prime_3_68 => 
            next_state <= square_with_reduction_special_prime_3_68;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_69;
            end if;
        when square_with_reduction_special_prime_3_69 => 
            next_state <= square_with_reduction_special_prime_3_69;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_70;
            end if;
        when square_with_reduction_special_prime_3_70 => 
            next_state <= square_with_reduction_special_prime_3_70;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_71;
            end if;
        when square_with_reduction_special_prime_3_71 => 
            next_state <= square_with_reduction_special_prime_3_71;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_72;
            end if;
        when square_with_reduction_special_prime_3_72 => 
            next_state <= square_with_reduction_special_prime_3_72;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_73;
            end if;
        when square_with_reduction_special_prime_3_73 => 
            next_state <= square_with_reduction_special_prime_3_73;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_74;
            end if;
        when square_with_reduction_special_prime_3_74 => 
            next_state <= square_with_reduction_special_prime_3_74;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_75;
            end if;
        when square_with_reduction_special_prime_3_75 => 
            next_state <= square_with_reduction_special_prime_3_75;
            if(ultimate_operation = '1') then
                if(operands_size = "110") then
                    next_state <= square_with_reduction_special_prime_3_76;
                else
                    next_state <= square_with_reduction_special_prime_3_108;
                end if;
            end if;
        when square_with_reduction_special_prime_3_76 => 
            next_state <= square_with_reduction_special_prime_3_76;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_77;
            end if;
        when square_with_reduction_special_prime_3_77 => 
            next_state <= square_with_reduction_special_prime_3_77;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_78;
            end if;
        when square_with_reduction_special_prime_3_78 => 
            next_state <= square_with_reduction_special_prime_3_78;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_79;
            end if;
        when square_with_reduction_special_prime_3_79 => 
            next_state <= square_with_reduction_special_prime_3_79;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_80;
            end if;
        when square_with_reduction_special_prime_3_80 => 
            next_state <= square_with_reduction_special_prime_3_80;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_81;
            end if;
        when square_with_reduction_special_prime_3_81 => 
            next_state <= square_with_reduction_special_prime_3_81;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_82;
            end if;
        when square_with_reduction_special_prime_3_82 => 
            next_state <= square_with_reduction_special_prime_3_82;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_83;
            end if;
        when square_with_reduction_special_prime_3_83 => 
            next_state <= square_with_reduction_special_prime_3_83;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_84;
            end if;
        when square_with_reduction_special_prime_3_84 => 
            next_state <= square_with_reduction_special_prime_3_84;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_85;
            end if;
        when square_with_reduction_special_prime_3_85 => 
            next_state <= square_with_reduction_special_prime_3_85;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_86;
            end if;
        when square_with_reduction_special_prime_3_86 => 
            next_state <= square_with_reduction_special_prime_3_86;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_87;
            end if;
        when square_with_reduction_special_prime_3_87 => 
            next_state <= square_with_reduction_special_prime_3_87;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_88;
            end if;
        when square_with_reduction_special_prime_3_88 => 
            next_state <= square_with_reduction_special_prime_3_88;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_89;
            end if;
        when square_with_reduction_special_prime_3_89 => 
            next_state <= square_with_reduction_special_prime_3_89;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_90;
            end if;
        when square_with_reduction_special_prime_3_90 => 
            next_state <= square_with_reduction_special_prime_3_90;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_91;
            end if;
        when square_with_reduction_special_prime_3_91 => 
            next_state <= square_with_reduction_special_prime_3_91;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_92;
            end if;
        when square_with_reduction_special_prime_3_92 => 
            next_state <= square_with_reduction_special_prime_3_92;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_93;
            end if;
        when square_with_reduction_special_prime_3_93 => 
            next_state <= square_with_reduction_special_prime_3_93;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_94;
            end if;
        when square_with_reduction_special_prime_3_94 => 
            next_state <= square_with_reduction_special_prime_3_94;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_95;
            end if;
        when square_with_reduction_special_prime_3_95 => 
            next_state <= square_with_reduction_special_prime_3_95;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_96;
            end if;
        when square_with_reduction_special_prime_3_96 => 
            next_state <= square_with_reduction_special_prime_3_96;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_97;
            end if;
        when square_with_reduction_special_prime_3_97 => 
            next_state <= square_with_reduction_special_prime_3_97;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_98;
            end if;
        when square_with_reduction_special_prime_3_98 => 
            next_state <= square_with_reduction_special_prime_3_98;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_99;
            end if;
        when square_with_reduction_special_prime_3_99 => 
            next_state <= square_with_reduction_special_prime_3_99;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_100;
            end if;
        when square_with_reduction_special_prime_3_100 => 
            next_state <= square_with_reduction_special_prime_3_100;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_101;
            end if;
        when square_with_reduction_special_prime_3_101 => 
            next_state <= square_with_reduction_special_prime_3_101;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_102;
            end if;
        when square_with_reduction_special_prime_3_102 => 
            next_state <= square_with_reduction_special_prime_3_102;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_103;
            end if;
        when square_with_reduction_special_prime_3_103 => 
            next_state <= square_with_reduction_special_prime_3_103;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_104;
            end if;
        when square_with_reduction_special_prime_3_104 => 
            next_state <= square_with_reduction_special_prime_3_104;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_105;
            end if;
        when square_with_reduction_special_prime_3_105 => 
            next_state <= square_with_reduction_special_prime_3_105;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_106;
            end if;            
        when square_with_reduction_special_prime_3_106 => 
            next_state <= square_with_reduction_special_prime_3_106;
            if(ultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when square_with_reduction_special_prime_3_108 => 
            next_state <= square_with_reduction_special_prime_3_108;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_109;
            end if;
        when square_with_reduction_special_prime_3_109 => 
            next_state <= square_with_reduction_special_prime_3_109;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_110;
            end if;
        when square_with_reduction_special_prime_3_110 => 
            next_state <= square_with_reduction_special_prime_3_110;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_111;
            end if;
        when square_with_reduction_special_prime_3_111 => 
            next_state <= square_with_reduction_special_prime_3_111;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_112;
            end if;
        when square_with_reduction_special_prime_3_112 => 
            next_state <= square_with_reduction_special_prime_3_112;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_113;
            end if;
        when square_with_reduction_special_prime_3_113 => 
            next_state <= square_with_reduction_special_prime_3_113;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_114;
            end if;
        when square_with_reduction_special_prime_3_114 => 
            next_state <= square_with_reduction_special_prime_3_114;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_115;
            end if;
        when square_with_reduction_special_prime_3_115 => 
            next_state <= square_with_reduction_special_prime_3_115;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_116;
            end if;
        when square_with_reduction_special_prime_3_116 => 
            next_state <= square_with_reduction_special_prime_3_116;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_117;
            end if;
        when square_with_reduction_special_prime_3_117 => 
            next_state <= square_with_reduction_special_prime_3_117;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_118;
            end if;
        when square_with_reduction_special_prime_3_118 => 
            next_state <= square_with_reduction_special_prime_3_118;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_119;
            end if;
        when square_with_reduction_special_prime_3_119 => 
            next_state <= square_with_reduction_special_prime_3_119;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_120;
            end if;
        when square_with_reduction_special_prime_3_120 => 
            next_state <= square_with_reduction_special_prime_3_120;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_121;
            end if;
        when square_with_reduction_special_prime_3_121 => 
            next_state <= square_with_reduction_special_prime_3_121;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_122;
            end if;
        when square_with_reduction_special_prime_3_122 => 
            next_state <= square_with_reduction_special_prime_3_122;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_123;
            end if;
        when square_with_reduction_special_prime_3_123 => 
            next_state <= square_with_reduction_special_prime_3_123;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_124;
            end if;
        when square_with_reduction_special_prime_3_124 => 
            next_state <= square_with_reduction_special_prime_3_124;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_125;
            end if;
        when square_with_reduction_special_prime_3_125 => 
            next_state <= square_with_reduction_special_prime_3_125;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_126;
            end if;
        when square_with_reduction_special_prime_3_126 => 
            next_state <= square_with_reduction_special_prime_3_126;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_127;
            end if;
        when square_with_reduction_special_prime_3_127 => 
            next_state <= square_with_reduction_special_prime_3_127;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_128;
            end if;
        when square_with_reduction_special_prime_3_128 => 
            next_state <= square_with_reduction_special_prime_3_128;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_129;
            end if;
        when square_with_reduction_special_prime_3_129 => 
            next_state <= square_with_reduction_special_prime_3_129;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_130;
            end if;
        when square_with_reduction_special_prime_3_130 => 
            next_state <= square_with_reduction_special_prime_3_130;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_131;
            end if;
        when square_with_reduction_special_prime_3_131 => 
            next_state <= square_with_reduction_special_prime_3_131;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_132;
            end if;
        when square_with_reduction_special_prime_3_132 => 
            next_state <= square_with_reduction_special_prime_3_132;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_133;
            end if;
        when square_with_reduction_special_prime_3_133 => 
            next_state <= square_with_reduction_special_prime_3_133;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_134;
            end if;
        when square_with_reduction_special_prime_3_134 => 
            next_state <= square_with_reduction_special_prime_3_134;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_135;
            end if;
        when square_with_reduction_special_prime_3_135 => 
            next_state <= square_with_reduction_special_prime_3_135;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_136;
            end if;
        when square_with_reduction_special_prime_3_136 => 
            next_state <= square_with_reduction_special_prime_3_136;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_137;
            end if;
        when square_with_reduction_special_prime_3_137 => 
            next_state <= square_with_reduction_special_prime_3_137;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_138;
            end if;
        when square_with_reduction_special_prime_3_138 => 
            next_state <= square_with_reduction_special_prime_3_138;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_139;
            end if;
        when square_with_reduction_special_prime_3_139 => 
            next_state <= square_with_reduction_special_prime_3_139;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_140;
            end if;
        when square_with_reduction_special_prime_3_140 => 
            next_state <= square_with_reduction_special_prime_3_140;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_141;
            end if;
        when square_with_reduction_special_prime_3_141 => 
            next_state <= square_with_reduction_special_prime_3_141;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_142;
            end if;
        when square_with_reduction_special_prime_3_142 => 
            next_state <= square_with_reduction_special_prime_3_142;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_143;
            end if;
        when square_with_reduction_special_prime_3_143 => 
            next_state <= square_with_reduction_special_prime_3_143;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_144;
            end if;
        when square_with_reduction_special_prime_3_144 => 
            next_state <= square_with_reduction_special_prime_3_144;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_145;
            end if;
        when square_with_reduction_special_prime_3_145 => 
            next_state <= square_with_reduction_special_prime_3_145;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_146;
            end if;
        when square_with_reduction_special_prime_3_146 => 
            next_state <= square_with_reduction_special_prime_3_146;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_147;
            end if;
        when square_with_reduction_special_prime_3_147 => 
            next_state <= square_with_reduction_special_prime_3_147;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_148;
            end if;
        when square_with_reduction_special_prime_3_148 => 
            next_state <= square_with_reduction_special_prime_3_148;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_149;
            end if;
        when square_with_reduction_special_prime_3_149 => 
            next_state <= square_with_reduction_special_prime_3_149;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_150;
            end if;
        when square_with_reduction_special_prime_3_150 => 
            next_state <= square_with_reduction_special_prime_3_150;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_151;
            end if;
        when square_with_reduction_special_prime_3_151 => 
            next_state <= square_with_reduction_special_prime_3_151;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_152;
            end if;
        when square_with_reduction_special_prime_3_152 => 
            next_state <= square_with_reduction_special_prime_3_152;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_153;
            end if;
        when square_with_reduction_special_prime_3_153 => 
            next_state <= square_with_reduction_special_prime_3_153;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_154;
            end if;
        when square_with_reduction_special_prime_3_154 => 
            next_state <= square_with_reduction_special_prime_3_154;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_155;
            end if;
        when square_with_reduction_special_prime_3_155 => 
            next_state <= square_with_reduction_special_prime_3_155;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_156;
            end if;
        when square_with_reduction_special_prime_3_156 => 
            next_state <= square_with_reduction_special_prime_3_156;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_157;
            end if;
        when square_with_reduction_special_prime_3_157 => 
            next_state <= square_with_reduction_special_prime_3_157;
            if(ultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_3_158;
            end if;
        when square_with_reduction_special_prime_3_158 => 
            next_state <= square_with_reduction_special_prime_3_158;
            if(ultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when addition_subtraction_direct_0 =>
            next_state <= addition_subtraction_direct_0;
            if(ultimate_operation = '1') then
                next_state <= nop_4_stages;
            end if;
        when addition_subtraction_direct_2 =>
            next_state <= addition_subtraction_direct_2;
            if(ultimate_operation = '1') then
                if(operands_size = "001") then
                    next_state <= addition_subtraction_direct_3;
                else
                    next_state <= addition_subtraction_direct_5;
                end if;
            end if;
        when addition_subtraction_direct_3 =>
            next_state <= addition_subtraction_direct_3;
            if(ultimate_operation = '1') then
                next_state <= nop_4_stages;
            end if;
        when addition_subtraction_direct_5 =>
            next_state <= addition_subtraction_direct_5;
            if(ultimate_operation = '1') then
                if(operands_size = "010") then
                    next_state <= addition_subtraction_direct_6;
                else
                    next_state <= addition_subtraction_direct_8;
                end if;
            end if;
        when addition_subtraction_direct_6 =>
            next_state <= addition_subtraction_direct_6;
            if(ultimate_operation = '1') then
                next_state <= nop_4_stages;
            end if;
        when addition_subtraction_direct_8 =>
            next_state <= addition_subtraction_direct_8;
            if(ultimate_operation = '1') then
                if(operands_size = "011") then
                    next_state <= addition_subtraction_direct_9;
                else
                    next_state <= addition_subtraction_direct_11;
                end if;
            end if;
        when addition_subtraction_direct_9 =>
            next_state <= addition_subtraction_direct_9;
            if(ultimate_operation = '1') then
                next_state <= nop_4_stages;
            end if;
        when addition_subtraction_direct_11 =>
            next_state <= addition_subtraction_direct_11;
            if(ultimate_operation = '1') then
                if(operands_size = "100") then
                    next_state <= addition_subtraction_direct_12;
                else
                    next_state <= addition_subtraction_direct_14;
                end if;
            end if;
        when addition_subtraction_direct_12 =>
            next_state <= addition_subtraction_direct_12;
            if(ultimate_operation = '1') then
                next_state <= nop_4_stages;
            end if;
        when addition_subtraction_direct_14 =>
            next_state <= addition_subtraction_direct_14;
            if(ultimate_operation = '1') then
                if(operands_size = "101") then
                    next_state <= addition_subtraction_direct_15;
                else
                    next_state <= addition_subtraction_direct_17;
                end if;
            end if;
        when addition_subtraction_direct_15 =>
            next_state <= addition_subtraction_direct_15;
            if(ultimate_operation = '1') then
                next_state <= nop_4_stages;
            end if;
        when addition_subtraction_direct_17 =>
            next_state <= addition_subtraction_direct_17;
            if(ultimate_operation = '1') then
                if(operands_size = "110") then
                    next_state <= addition_subtraction_direct_18;
                else
                    next_state <= addition_subtraction_direct_20;
                end if;
            end if;
        when addition_subtraction_direct_18 =>
            next_state <= addition_subtraction_direct_18;
            if(ultimate_operation = '1') then
                next_state <= nop_4_stages;
            end if;
        when addition_subtraction_direct_20 =>
            next_state <= addition_subtraction_direct_20;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_direct_21;
            end if;
        when addition_subtraction_direct_21 =>
            next_state <= addition_subtraction_direct_21;
            if(ultimate_operation = '1') then
                next_state <= nop_4_stages;
            end if;
        when iterative_modular_reduction_0 =>
            next_state <= iterative_modular_reduction_0;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_1;
            end if;    
        when iterative_modular_reduction_1 =>
            next_state <= iterative_modular_reduction_1;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_2;
            end if;
        when iterative_modular_reduction_2 =>
            next_state <= iterative_modular_reduction_2;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_3;
            end if;
        when iterative_modular_reduction_3 =>
            next_state <= iterative_modular_reduction_3;
            if(ultimate_operation = '1') then
                next_state <= nop_4_stages;
            end if;
        when iterative_modular_reduction_5 =>
            next_state <= iterative_modular_reduction_5;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_6;
            end if;
        when iterative_modular_reduction_6 =>
            next_state <= iterative_modular_reduction_6;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_7;
            end if;
        when iterative_modular_reduction_7 =>
            next_state <= iterative_modular_reduction_7;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_8;
            end if;
        when iterative_modular_reduction_8 =>
            next_state <= iterative_modular_reduction_8;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_9;
            end if;
        when iterative_modular_reduction_9 =>
            next_state <= iterative_modular_reduction_9;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_10;
            end if;
        when iterative_modular_reduction_10 =>
            next_state <= iterative_modular_reduction_10;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_11;
            end if;
        when iterative_modular_reduction_11 =>
            next_state <= iterative_modular_reduction_11;
            if(ultimate_operation = '1') then
                next_state <= nop_4_stages;
            end if;
        when iterative_modular_reduction_13 =>
            next_state <= iterative_modular_reduction_13;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_14;
            end if;
        when iterative_modular_reduction_14 =>
            next_state <= iterative_modular_reduction_14;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_15;
            end if;
        when iterative_modular_reduction_15 =>
            next_state <= iterative_modular_reduction_15;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_16;
            end if;
        when iterative_modular_reduction_16 =>
            next_state <= iterative_modular_reduction_16;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_17;
            end if;
        when iterative_modular_reduction_17 =>
            next_state <= iterative_modular_reduction_17;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_18;
            end if;
        when iterative_modular_reduction_18 =>
            next_state <= iterative_modular_reduction_18;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_19;
            end if;
        when iterative_modular_reduction_19 =>
            next_state <= iterative_modular_reduction_19;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_20;
            end if;
        when iterative_modular_reduction_20 =>
            next_state <= iterative_modular_reduction_20;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_21;
            end if;
        when iterative_modular_reduction_21 =>
            next_state <= iterative_modular_reduction_21;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_22;
            end if;
        when iterative_modular_reduction_22 =>
            next_state <= iterative_modular_reduction_22;
            if(ultimate_operation = '1') then
                next_state <= nop_4_stages;
            end if;
        when iterative_modular_reduction_24 =>
            next_state <= iterative_modular_reduction_24;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_25;
            end if;
        when iterative_modular_reduction_25 =>
            next_state <= iterative_modular_reduction_25;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_26;
            end if;
        when iterative_modular_reduction_26 =>
            next_state <= iterative_modular_reduction_26;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_27;
            end if;
        when iterative_modular_reduction_27 =>
            next_state <= iterative_modular_reduction_27;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_28;
            end if;
        when iterative_modular_reduction_28 =>
            next_state <= iterative_modular_reduction_28;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_29;
            end if;
        when iterative_modular_reduction_29 =>
            next_state <= iterative_modular_reduction_29;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_30;
            end if;
        when iterative_modular_reduction_30 =>
            next_state <= iterative_modular_reduction_30;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_31;
            end if;
        when iterative_modular_reduction_31 =>
            next_state <= iterative_modular_reduction_31;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_32;
            end if;
        when iterative_modular_reduction_32 =>
            next_state <= iterative_modular_reduction_32;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_33;
            end if;
        when iterative_modular_reduction_33 =>
            next_state <= iterative_modular_reduction_33;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_34;
            end if;
        when iterative_modular_reduction_34 =>
            next_state <= iterative_modular_reduction_34;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_35;
            end if;
        when iterative_modular_reduction_35 =>
            next_state <= iterative_modular_reduction_35;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_36;
            end if;
        when iterative_modular_reduction_36 =>
            next_state <= iterative_modular_reduction_36;
            if(ultimate_operation = '1') then
                next_state <= nop_4_stages;
            end if;
        when iterative_modular_reduction_38 =>
            next_state <= iterative_modular_reduction_38;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_39;
            end if;
        when iterative_modular_reduction_39 =>
            next_state <= iterative_modular_reduction_39;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_40;
            end if;
        when iterative_modular_reduction_40 =>
            next_state <= iterative_modular_reduction_40;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_41;
            end if;
        when iterative_modular_reduction_41 =>
            next_state <= iterative_modular_reduction_41;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_42;
            end if;
        when iterative_modular_reduction_42 =>
            next_state <= iterative_modular_reduction_42;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_43;
            end if;
        when iterative_modular_reduction_43 =>
            next_state <= iterative_modular_reduction_43;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_44;
            end if;
        when iterative_modular_reduction_44 =>
            next_state <= iterative_modular_reduction_44;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_45;
            end if;
        when iterative_modular_reduction_45 =>
            next_state <= iterative_modular_reduction_45;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_46;
            end if;
        when iterative_modular_reduction_46 =>
            next_state <= iterative_modular_reduction_46;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_47;
            end if;
        when iterative_modular_reduction_47 =>
            next_state <= iterative_modular_reduction_47;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_48;
            end if;
        when iterative_modular_reduction_48 =>
            next_state <= iterative_modular_reduction_48;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_49;
            end if;
        when iterative_modular_reduction_49 =>
            next_state <= iterative_modular_reduction_49;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_50;
            end if;
        when iterative_modular_reduction_50 =>
            next_state <= iterative_modular_reduction_50;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_51;
            end if;
        when iterative_modular_reduction_51 =>
            next_state <= iterative_modular_reduction_51;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_52;
            end if;
        when iterative_modular_reduction_52 =>
            next_state <= iterative_modular_reduction_52;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_53;
            end if;
        when iterative_modular_reduction_53 =>
            next_state <= iterative_modular_reduction_53;
            if(ultimate_operation = '1') then
                next_state <= nop_4_stages;
            end if;
        when iterative_modular_reduction_55 =>
            next_state <= iterative_modular_reduction_55;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_56;
            end if;
        when iterative_modular_reduction_56 =>
            next_state <= iterative_modular_reduction_56;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_57;
            end if;
        when iterative_modular_reduction_57 =>
            next_state <= iterative_modular_reduction_57;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_58;
            end if;
        when iterative_modular_reduction_58 =>
            next_state <= iterative_modular_reduction_58;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_59;
            end if;
        when iterative_modular_reduction_59 =>
            next_state <= iterative_modular_reduction_59;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_60;
            end if;
        when iterative_modular_reduction_60 =>
            next_state <= iterative_modular_reduction_60;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_61;
            end if;
        when iterative_modular_reduction_61 =>
            next_state <= iterative_modular_reduction_61;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_62;
            end if;
        when iterative_modular_reduction_62 =>
            next_state <= iterative_modular_reduction_62;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_63;
            end if;
        when iterative_modular_reduction_63 =>
            next_state <= iterative_modular_reduction_63;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_64;
            end if;
        when iterative_modular_reduction_64 =>
            next_state <= iterative_modular_reduction_64;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_65;
            end if;
        when iterative_modular_reduction_65 =>
            next_state <= iterative_modular_reduction_65;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_66;
            end if;
        when iterative_modular_reduction_66 =>
            next_state <= iterative_modular_reduction_66;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_67;
            end if;
        when iterative_modular_reduction_67 =>
            next_state <= iterative_modular_reduction_67;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_68;
            end if;
        when iterative_modular_reduction_68 =>
            next_state <= iterative_modular_reduction_68;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_69;
            end if;
        when iterative_modular_reduction_69 =>
            next_state <= iterative_modular_reduction_69;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_70;
            end if;
        when iterative_modular_reduction_70 =>
            next_state <= iterative_modular_reduction_70;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_71;
            end if;
        when iterative_modular_reduction_71 =>
            next_state <= iterative_modular_reduction_71;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_72;
            end if;
        when iterative_modular_reduction_72 =>
            next_state <= iterative_modular_reduction_72;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_73;
            end if;
        when iterative_modular_reduction_73 =>
            next_state <= iterative_modular_reduction_73;
            if(ultimate_operation = '1') then
                next_state <= nop_4_stages;
            end if;
        when iterative_modular_reduction_75 =>
            next_state <= iterative_modular_reduction_75;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_76;
            end if;
        when iterative_modular_reduction_76 =>
            next_state <= iterative_modular_reduction_76;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_77;
            end if;
        when iterative_modular_reduction_77 =>
            next_state <= iterative_modular_reduction_77;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_78;
            end if;
        when iterative_modular_reduction_78 =>
            next_state <= iterative_modular_reduction_78;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_79;
            end if;
        when iterative_modular_reduction_79 =>
            next_state <= iterative_modular_reduction_79;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_80;
            end if;
        when iterative_modular_reduction_80 =>
            next_state <= iterative_modular_reduction_80;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_81;
            end if;
        when iterative_modular_reduction_81 =>
            next_state <= iterative_modular_reduction_81;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_82;
            end if;
        when iterative_modular_reduction_82 =>
            next_state <= iterative_modular_reduction_82;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_83;
            end if;
        when iterative_modular_reduction_83 =>
            next_state <= iterative_modular_reduction_83;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_84;
            end if;
        when iterative_modular_reduction_84 =>
            next_state <= iterative_modular_reduction_84;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_85;
            end if;
        when iterative_modular_reduction_85 =>
            next_state <= iterative_modular_reduction_85;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_86;
            end if;
        when iterative_modular_reduction_86 =>
            next_state <= iterative_modular_reduction_86;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_87;
            end if;
        when iterative_modular_reduction_87 =>
            next_state <= iterative_modular_reduction_87;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_88;
            end if;
        when iterative_modular_reduction_88 =>
            next_state <= iterative_modular_reduction_88;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_89;
            end if;
        when iterative_modular_reduction_89 =>
            next_state <= iterative_modular_reduction_89;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_90;
            end if;
        when iterative_modular_reduction_90 =>
            next_state <= iterative_modular_reduction_90;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_91;
            end if;
        when iterative_modular_reduction_91 =>
            next_state <= iterative_modular_reduction_91;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_92;
            end if;
        when iterative_modular_reduction_92 =>
            next_state <= iterative_modular_reduction_92;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_93;
            end if;
        when iterative_modular_reduction_93 =>
            next_state <= iterative_modular_reduction_93;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_94;
            end if;
        when iterative_modular_reduction_94 =>
            next_state <= iterative_modular_reduction_94;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_95;
            end if;
        when iterative_modular_reduction_95 =>
            next_state <= iterative_modular_reduction_95;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_96;
            end if;
        when iterative_modular_reduction_96 =>
            next_state <= iterative_modular_reduction_96;
            if(ultimate_operation = '1') then
                next_state <= nop_4_stages;
            end if;
        when iterative_modular_reduction_98 =>
            next_state <= iterative_modular_reduction_98;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_99;
            end if;
        when iterative_modular_reduction_99 =>
            next_state <= iterative_modular_reduction_99;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_100;
            end if;
        when iterative_modular_reduction_100 =>
            next_state <= iterative_modular_reduction_100;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_101;
            end if;
        when iterative_modular_reduction_101 =>
            next_state <= iterative_modular_reduction_101;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_102;
            end if;
        when iterative_modular_reduction_102 =>
            next_state <= iterative_modular_reduction_102;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_103;
            end if;
        when iterative_modular_reduction_103 =>
            next_state <= iterative_modular_reduction_103;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_104;
            end if;
        when iterative_modular_reduction_104 =>
            next_state <= iterative_modular_reduction_104;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_105;
            end if;
        when iterative_modular_reduction_105 =>
            next_state <= iterative_modular_reduction_105;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_106;
            end if;
        when iterative_modular_reduction_106 =>
            next_state <= iterative_modular_reduction_106;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_107;
            end if;
        when iterative_modular_reduction_107 =>
            next_state <= iterative_modular_reduction_107;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_108;
            end if;
        when iterative_modular_reduction_108 =>
            next_state <= iterative_modular_reduction_108;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_109;
            end if;
        when iterative_modular_reduction_109 =>
            next_state <= iterative_modular_reduction_109;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_110;
            end if;
        when iterative_modular_reduction_110 =>
            next_state <= iterative_modular_reduction_110;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_111;
            end if;
        when iterative_modular_reduction_111 =>
            next_state <= iterative_modular_reduction_111;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_112;
            end if;
        when iterative_modular_reduction_112 =>
            next_state <= iterative_modular_reduction_112;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_113;
            end if;
        when iterative_modular_reduction_113 =>
            next_state <= iterative_modular_reduction_113;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_114;
            end if;
        when iterative_modular_reduction_114 =>
            next_state <= iterative_modular_reduction_114;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_115;
            end if;
        when iterative_modular_reduction_115 =>
            next_state <= iterative_modular_reduction_115;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_116;
            end if;
        when iterative_modular_reduction_116 =>
            next_state <= iterative_modular_reduction_116;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_117;
            end if;
        when iterative_modular_reduction_117 =>
            next_state <= iterative_modular_reduction_117;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_118;
            end if;
        when iterative_modular_reduction_118 =>
            next_state <= iterative_modular_reduction_118;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_119;
            end if;
        when iterative_modular_reduction_119 =>
            next_state <= iterative_modular_reduction_119;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_120;
            end if;
        when iterative_modular_reduction_120 =>
            next_state <= iterative_modular_reduction_120;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_121;
            end if;
        when iterative_modular_reduction_121 =>
            next_state <= iterative_modular_reduction_121;
            if(ultimate_operation = '1') then
                next_state <= iterative_modular_reduction_122;
            end if;
        when iterative_modular_reduction_122 =>
            next_state <= iterative_modular_reduction_122;
            if(ultimate_operation = '1') then
                next_state <= nop_4_stages;
            end if;
        when addition_subtraction_with_reduction_0 =>
            next_state <= addition_subtraction_with_reduction_0;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_1;
            end if;
        when addition_subtraction_with_reduction_1 =>
            next_state <= addition_subtraction_with_reduction_1;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_2;
            end if;
        when addition_subtraction_with_reduction_2 =>
            next_state <= addition_subtraction_with_reduction_2;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_3;
            end if;
        when addition_subtraction_with_reduction_3 =>
            next_state <= addition_subtraction_with_reduction_3;
            if(ultimate_operation = '1') then
                next_state <= nop_4_stages;
            end if;
        when addition_subtraction_with_reduction_5 =>
            next_state <= addition_subtraction_with_reduction_5;
            if(ultimate_operation = '1') then
                if(operands_size = "001") then
                    next_state <= addition_subtraction_with_reduction_6;
                else
                    next_state <= addition_subtraction_with_reduction_14;
                end if;
            end if;
        when addition_subtraction_with_reduction_6 =>
            next_state <= addition_subtraction_with_reduction_6;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_7;
            end if;
        when addition_subtraction_with_reduction_7 =>
            next_state <= addition_subtraction_with_reduction_7;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_8;
            end if;
        when addition_subtraction_with_reduction_8 =>
            next_state <= addition_subtraction_with_reduction_8;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_9;
            end if;
        when addition_subtraction_with_reduction_9 =>
            next_state <= addition_subtraction_with_reduction_9;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_10;
            end if;
        when addition_subtraction_with_reduction_10 =>
            next_state <= addition_subtraction_with_reduction_10;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_11;
            end if;
        when addition_subtraction_with_reduction_11 =>
            next_state <= addition_subtraction_with_reduction_11;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_12;
            end if;
        when addition_subtraction_with_reduction_12 =>
            next_state <= addition_subtraction_with_reduction_12;
            if(ultimate_operation = '1') then
                next_state <= nop_4_stages;
            end if;
        when addition_subtraction_with_reduction_14 =>
            next_state <= addition_subtraction_with_reduction_14;
            if(ultimate_operation = '1') then
                if(operands_size = "010") then
                    next_state <= addition_subtraction_with_reduction_15;
                else
                    next_state <= addition_subtraction_with_reduction_26;
                end if;
            end if;
        when addition_subtraction_with_reduction_15 =>
            next_state <= addition_subtraction_with_reduction_15;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_16;
            end if;
        when addition_subtraction_with_reduction_16 =>
            next_state <= addition_subtraction_with_reduction_16;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_17;
            end if;
        when addition_subtraction_with_reduction_17 =>
            next_state <= addition_subtraction_with_reduction_17;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_18;
            end if;
        when addition_subtraction_with_reduction_18 =>
            next_state <= addition_subtraction_with_reduction_18;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_19;
            end if;
        when addition_subtraction_with_reduction_19 =>
            next_state <= addition_subtraction_with_reduction_19;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_20;
            end if;
        when addition_subtraction_with_reduction_20 =>
            next_state <= addition_subtraction_with_reduction_20;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_21;
            end if;
        when addition_subtraction_with_reduction_21 =>
            next_state <= addition_subtraction_with_reduction_21;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_22;
            end if;
        when addition_subtraction_with_reduction_22 =>
            next_state <= addition_subtraction_with_reduction_22;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_23;
            end if;
        when addition_subtraction_with_reduction_23 =>
            next_state <= addition_subtraction_with_reduction_23;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_24;
            end if;
        when addition_subtraction_with_reduction_24 =>
            next_state <= addition_subtraction_with_reduction_24;
            if(ultimate_operation = '1') then
                next_state <= nop_4_stages;
            end if;
        when addition_subtraction_with_reduction_26 =>
            next_state <= addition_subtraction_with_reduction_26;
            if(ultimate_operation = '1') then
                if(operands_size = "011") then
                    next_state <= addition_subtraction_with_reduction_27;
                else
                    next_state <= addition_subtraction_with_reduction_41;
                end if;
            end if;
        when addition_subtraction_with_reduction_27 =>
            next_state <= addition_subtraction_with_reduction_27;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_28;
            end if;
        when addition_subtraction_with_reduction_28 =>
            next_state <= addition_subtraction_with_reduction_28;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_29;
            end if;
        when addition_subtraction_with_reduction_29 =>
            next_state <= addition_subtraction_with_reduction_29;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_30;
            end if;
        when addition_subtraction_with_reduction_30 =>
            next_state <= addition_subtraction_with_reduction_30;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_31;
            end if;
        when addition_subtraction_with_reduction_31 =>
            next_state <= addition_subtraction_with_reduction_31;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_32;
            end if;
        when addition_subtraction_with_reduction_32 =>
            next_state <= addition_subtraction_with_reduction_32;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_33;
            end if;
        when addition_subtraction_with_reduction_33 =>
            next_state <= addition_subtraction_with_reduction_33;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_34;
            end if;
        when addition_subtraction_with_reduction_34 =>
            next_state <= addition_subtraction_with_reduction_34;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_35;
            end if;
        when addition_subtraction_with_reduction_35 =>
            next_state <= addition_subtraction_with_reduction_35;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_36;
            end if;
        when addition_subtraction_with_reduction_36 =>
            next_state <= addition_subtraction_with_reduction_36;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_37;
            end if;
        when addition_subtraction_with_reduction_37 =>
            next_state <= addition_subtraction_with_reduction_37;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_38;
            end if;
        when addition_subtraction_with_reduction_38 =>
            next_state <= addition_subtraction_with_reduction_38;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_39;
            end if;
        when addition_subtraction_with_reduction_39 =>
            next_state <= addition_subtraction_with_reduction_39;
            if(ultimate_operation = '1') then
                next_state <= nop_4_stages;
            end if;
        when addition_subtraction_with_reduction_41 =>
            next_state <= addition_subtraction_with_reduction_41;
            if(ultimate_operation = '1') then
                if(operands_size = "100") then
                    next_state <= addition_subtraction_with_reduction_42;
                else
                    next_state <= addition_subtraction_with_reduction_59;
                end if;
            end if;
        when addition_subtraction_with_reduction_42 =>
            next_state <= addition_subtraction_with_reduction_42;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_43;
            end if;
        when addition_subtraction_with_reduction_43 =>
            next_state <= addition_subtraction_with_reduction_43;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_44;
            end if;
        when addition_subtraction_with_reduction_44 =>
            next_state <= addition_subtraction_with_reduction_44;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_45;
            end if;
        when addition_subtraction_with_reduction_45 =>
            next_state <= addition_subtraction_with_reduction_45;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_46;
            end if;
        when addition_subtraction_with_reduction_46 =>
            next_state <= addition_subtraction_with_reduction_46;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_47;
            end if;
        when addition_subtraction_with_reduction_47 =>
            next_state <= addition_subtraction_with_reduction_47;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_48;
            end if;
        when addition_subtraction_with_reduction_48 =>
            next_state <= addition_subtraction_with_reduction_48;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_49;
            end if;
        when addition_subtraction_with_reduction_49 =>
            next_state <= addition_subtraction_with_reduction_49;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_50;
            end if;
        when addition_subtraction_with_reduction_50 =>
            next_state <= addition_subtraction_with_reduction_50;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_51;
            end if;
        when addition_subtraction_with_reduction_51 =>
            next_state <= addition_subtraction_with_reduction_51;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_52;
            end if;
        when addition_subtraction_with_reduction_52 =>
            next_state <= addition_subtraction_with_reduction_52;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_53;
            end if;
        when addition_subtraction_with_reduction_53 =>
            next_state <= addition_subtraction_with_reduction_53;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_54;
            end if;
        when addition_subtraction_with_reduction_54 =>
            next_state <= addition_subtraction_with_reduction_54;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_55;
            end if;
        when addition_subtraction_with_reduction_55 =>
            next_state <= addition_subtraction_with_reduction_55;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_56;
            end if;
        when addition_subtraction_with_reduction_56 =>
            next_state <= addition_subtraction_with_reduction_56;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_57;
            end if;
        when addition_subtraction_with_reduction_57 =>
            next_state <= addition_subtraction_with_reduction_57;
            if(ultimate_operation = '1') then
                next_state <= nop_4_stages;
            end if;
        when addition_subtraction_with_reduction_59 =>
            next_state <= addition_subtraction_with_reduction_59;
            if(ultimate_operation = '1') then
                if(operands_size = "101") then
                    next_state <= addition_subtraction_with_reduction_60;
                else
                    next_state <= addition_subtraction_with_reduction_80;
                end if;
            end if;
        when addition_subtraction_with_reduction_60 =>
            next_state <= addition_subtraction_with_reduction_60;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_61;
            end if;
        when addition_subtraction_with_reduction_61 =>
            next_state <= addition_subtraction_with_reduction_61;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_62;
            end if;
        when addition_subtraction_with_reduction_62 =>
            next_state <= addition_subtraction_with_reduction_62;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_63;
            end if;
        when addition_subtraction_with_reduction_63 =>
            next_state <= addition_subtraction_with_reduction_63;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_64;
            end if;
        when addition_subtraction_with_reduction_64 =>
            next_state <= addition_subtraction_with_reduction_64;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_65;
            end if;
        when addition_subtraction_with_reduction_65 =>
            next_state <= addition_subtraction_with_reduction_65;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_66;
            end if;
        when addition_subtraction_with_reduction_66 =>
            next_state <= addition_subtraction_with_reduction_66;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_67;
            end if;
        when addition_subtraction_with_reduction_67 =>
            next_state <= addition_subtraction_with_reduction_67;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_68;
            end if;
        when addition_subtraction_with_reduction_68 =>
            next_state <= addition_subtraction_with_reduction_68;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_69;
            end if;
        when addition_subtraction_with_reduction_69 =>
            next_state <= addition_subtraction_with_reduction_69;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_70;
            end if;
        when addition_subtraction_with_reduction_70 =>
            next_state <= addition_subtraction_with_reduction_70;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_71;
            end if;
        when addition_subtraction_with_reduction_71 =>
            next_state <= addition_subtraction_with_reduction_71;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_72;
            end if;
        when addition_subtraction_with_reduction_72 =>
            next_state <= addition_subtraction_with_reduction_72;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_73;
            end if;
        when addition_subtraction_with_reduction_73 =>
            next_state <= addition_subtraction_with_reduction_73;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_74;
            end if;
        when addition_subtraction_with_reduction_74 =>
            next_state <= addition_subtraction_with_reduction_74;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_75;
            end if;
        when addition_subtraction_with_reduction_75 =>
            next_state <= addition_subtraction_with_reduction_75;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_76;
            end if;
        when addition_subtraction_with_reduction_76 =>
            next_state <= addition_subtraction_with_reduction_76;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_77;
            end if;
        when addition_subtraction_with_reduction_77 =>
            next_state <= addition_subtraction_with_reduction_77;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_78;
            end if;
        when addition_subtraction_with_reduction_78 =>
            next_state <= addition_subtraction_with_reduction_78;
            if(ultimate_operation = '1') then
                next_state <= nop_4_stages;
            end if;
        when addition_subtraction_with_reduction_80 =>
            next_state <= addition_subtraction_with_reduction_80;
            if(ultimate_operation = '1') then
                if(operands_size = "110") then
                    next_state <= addition_subtraction_with_reduction_81;
                else
                    next_state <= addition_subtraction_with_reduction_104;
                end if;
            end if;
        when addition_subtraction_with_reduction_81 =>
            next_state <= addition_subtraction_with_reduction_81;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_82;
            end if;
        when addition_subtraction_with_reduction_82 =>
            next_state <= addition_subtraction_with_reduction_82;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_83;
            end if;
        when addition_subtraction_with_reduction_83 =>
            next_state <= addition_subtraction_with_reduction_83;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_84;
            end if;
        when addition_subtraction_with_reduction_84 =>
            next_state <= addition_subtraction_with_reduction_84;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_85;
            end if;
        when addition_subtraction_with_reduction_85 =>
            next_state <= addition_subtraction_with_reduction_85;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_86;
            end if;
        when addition_subtraction_with_reduction_86 =>
            next_state <= addition_subtraction_with_reduction_86;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_87;
            end if;
        when addition_subtraction_with_reduction_87 =>
            next_state <= addition_subtraction_with_reduction_87;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_88;
            end if;
        when addition_subtraction_with_reduction_88 =>
            next_state <= addition_subtraction_with_reduction_88;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_89;
            end if;
        when addition_subtraction_with_reduction_89 =>
            next_state <= addition_subtraction_with_reduction_89;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_90;
            end if;
        when addition_subtraction_with_reduction_90 =>
            next_state <= addition_subtraction_with_reduction_90;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_91;
            end if;
        when addition_subtraction_with_reduction_91 =>
            next_state <= addition_subtraction_with_reduction_91;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_92;
            end if;
        when addition_subtraction_with_reduction_92 =>
            next_state <= addition_subtraction_with_reduction_92;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_93;
            end if;
        when addition_subtraction_with_reduction_93 =>
            next_state <= addition_subtraction_with_reduction_93;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_94;
            end if;
        when addition_subtraction_with_reduction_94 =>
            next_state <= addition_subtraction_with_reduction_94;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_95;
            end if;
        when addition_subtraction_with_reduction_95 =>
            next_state <= addition_subtraction_with_reduction_95;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_96;
            end if;
        when addition_subtraction_with_reduction_96 =>
            next_state <= addition_subtraction_with_reduction_96;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_97;
            end if;
        when addition_subtraction_with_reduction_97 =>
            next_state <= addition_subtraction_with_reduction_97;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_98;
            end if;
        when addition_subtraction_with_reduction_98 =>
            next_state <= addition_subtraction_with_reduction_98;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_99;
            end if;
        when addition_subtraction_with_reduction_99 =>
            next_state <= addition_subtraction_with_reduction_99;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_100;
            end if;
        when addition_subtraction_with_reduction_100 =>
            next_state <= addition_subtraction_with_reduction_100;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_101;
            end if;
        when addition_subtraction_with_reduction_101 =>
            next_state <= addition_subtraction_with_reduction_101;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_102;
            end if;
        when addition_subtraction_with_reduction_102 =>
            next_state <= addition_subtraction_with_reduction_102;
            if(ultimate_operation = '1') then
                next_state <= nop_4_stages;
            end if;
        when addition_subtraction_with_reduction_104 =>
            next_state <= addition_subtraction_with_reduction_104;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_105;
            end if;
        when addition_subtraction_with_reduction_105 =>
            next_state <= addition_subtraction_with_reduction_105;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_106;
            end if;
        when addition_subtraction_with_reduction_106 =>
            next_state <= addition_subtraction_with_reduction_106;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_107;
            end if;
        when addition_subtraction_with_reduction_107 =>
            next_state <= addition_subtraction_with_reduction_107;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_108;
            end if;
        when addition_subtraction_with_reduction_108 =>
            next_state <= addition_subtraction_with_reduction_108;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_109;
            end if;
        when addition_subtraction_with_reduction_109 =>
            next_state <= addition_subtraction_with_reduction_109;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_110;
            end if;
        when addition_subtraction_with_reduction_110 =>
            next_state <= addition_subtraction_with_reduction_110;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_111;
            end if;
        when addition_subtraction_with_reduction_111 =>
            next_state <= addition_subtraction_with_reduction_111;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_112;
            end if;
        when addition_subtraction_with_reduction_112 =>
            next_state <= addition_subtraction_with_reduction_112;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_113;
            end if;
        when addition_subtraction_with_reduction_113 =>
            next_state <= addition_subtraction_with_reduction_113;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_114;
            end if;
        when addition_subtraction_with_reduction_114 =>
            next_state <= addition_subtraction_with_reduction_114;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_115;
            end if;
        when addition_subtraction_with_reduction_115 =>
            next_state <= addition_subtraction_with_reduction_115;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_116;
            end if;
        when addition_subtraction_with_reduction_116 =>
            next_state <= addition_subtraction_with_reduction_116;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_117;
            end if;
        when addition_subtraction_with_reduction_117 =>
            next_state <= addition_subtraction_with_reduction_117;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_118;
            end if;
        when addition_subtraction_with_reduction_118 =>
            next_state <= addition_subtraction_with_reduction_118;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_119;
            end if;
        when addition_subtraction_with_reduction_119 =>
            next_state <= addition_subtraction_with_reduction_119;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_120;
            end if;
        when addition_subtraction_with_reduction_120 =>
            next_state <= addition_subtraction_with_reduction_120;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_121;
            end if;
        when addition_subtraction_with_reduction_121 =>
            next_state <= addition_subtraction_with_reduction_121;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_122;
            end if;
        when addition_subtraction_with_reduction_122 =>
            next_state <= addition_subtraction_with_reduction_122;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_123;
            end if;
        when addition_subtraction_with_reduction_123 =>
            next_state <= addition_subtraction_with_reduction_123;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_124;
            end if;
        when addition_subtraction_with_reduction_124 =>
            next_state <= addition_subtraction_with_reduction_124;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_125;
            end if;
        when addition_subtraction_with_reduction_125 =>
            next_state <= addition_subtraction_with_reduction_125;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_126;
            end if;
        when addition_subtraction_with_reduction_126 =>
            next_state <= addition_subtraction_with_reduction_126;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_127;
            end if;
        when addition_subtraction_with_reduction_127 =>
            next_state <= addition_subtraction_with_reduction_127;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_128;
            end if;
        when addition_subtraction_with_reduction_128 =>
            next_state <= addition_subtraction_with_reduction_128;
            if(ultimate_operation = '1') then
                next_state <= addition_subtraction_with_reduction_129;
            end if;
        when addition_subtraction_with_reduction_129 =>
            next_state <= addition_subtraction_with_reduction_129;
            if(ultimate_operation = '1') then
                next_state <= nop_4_stages;
            end if;
        when nop_4_stages =>
            next_state <= nop_4_stages;
            if(ultimate_operation = '1') then
                next_state <= decode_instruction;
            end if;
        when nop_8_stages =>
            next_state <= nop_8_stages;
            if(ultimate_operation = '1') then
                next_state <= decode_instruction;
            end if;
    end case;
end process;

end behavioral;