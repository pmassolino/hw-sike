--
-- Implementation by Pedro Maat C. Massolino, hereby denoted as "the implementer".
--
-- To the extent possible under law, the implementer has waived all copyright
-- and related or neighboring rights to the source code in this file.
-- http://creativecommons.org/publicdomain/zero/1.0/
--
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity carmela_state_machine_v128 is
    Port (
        clk : in std_logic;
        rstn : in std_logic;
        instruction_values_valid : in std_logic;
        instruction_type : in std_logic_vector(3 downto 0);
        operands_size : in std_logic_vector(2 downto 0);
        prime_line_equal_one : in std_logic;
        penultimate_operation : in std_logic;
        sm_rotation_size : out std_logic_vector(1 downto 0);
        sm_circular_shift_enable : out std_logic;
        sel_address_a : out std_logic;
        sel_address_b_prime : out std_logic_vector(1 downto 0);
        sm_specific_mac_address_a : out std_logic_vector(2 downto 0);
        sm_specific_mac_address_b : out std_logic_vector(2 downto 0);
        sm_specific_mac_address_o : out std_logic_vector(2 downto 0);
        sm_specific_mac_next_address_o : out std_logic_vector(2 downto 0);
        mac_enable_signed_a : out std_logic;
        mac_enable_signed_b : out std_logic;
        mac_sel_load_reg_a : out std_logic_vector(1 downto 0);
        mac_clear_reg_b : out std_logic;
        mac_clear_reg_acc : out std_logic;
        mac_sel_shift_reg_o : out std_logic;
        mac_enable_update_reg_s : out std_logic;
        mac_sel_reg_s_reg_o_sign : out std_logic;
        mac_reg_s_reg_o_positive : out std_logic;
        sm_sign_a_mode : out std_logic;
        sm_mac_operation_mode : out std_logic_vector(1 downto 0);
        mac_enable_reg_s_mask : out std_logic;
        mac_subtraction_reg_a_b : out std_logic;
        mac_sel_multiply_two_a_b : out std_logic;
        mac_sel_reg_y_output : out std_logic;
        sm_mac_write_enable_output : out std_logic;
        mac_memory_double_mode : out std_logic;
        mac_memory_only_write_mode : out std_logic;
        base_address_generator_o_increment_previous_address : out std_logic;
        sm_free_flag : out std_logic
    );
end carmela_state_machine_v128;

architecture behavioral of carmela_state_machine_v128 is

type state is (reset, decode_instruction,
-- 0000 multiplication with no reduction
multiplication_direct_0,
multiplication_direct_2, multiplication_direct_3, multiplication_direct_4, multiplication_direct_5,
multiplication_direct_7, multiplication_direct_8, multiplication_direct_9, multiplication_direct_10, multiplication_direct_11, multiplication_direct_12, multiplication_direct_13, multiplication_direct_14,
multiplication_direct_16, multiplication_direct_17, multiplication_direct_18, multiplication_direct_19, multiplication_direct_20, multiplication_direct_21, multiplication_direct_22, multiplication_direct_23, multiplication_direct_24, multiplication_direct_25, multiplication_direct_26, multiplication_direct_27,
multiplication_direct_29, multiplication_direct_30, multiplication_direct_31, multiplication_direct_32, multiplication_direct_33, multiplication_direct_34, multiplication_direct_35, multiplication_direct_36, multiplication_direct_37, multiplication_direct_38, multiplication_direct_39, multiplication_direct_40, multiplication_direct_41, multiplication_direct_42, multiplication_direct_43, multiplication_direct_44, multiplication_direct_45,
multiplication_direct_47, multiplication_direct_48, multiplication_direct_49, multiplication_direct_50, multiplication_direct_51, multiplication_direct_52, multiplication_direct_53, multiplication_direct_54, multiplication_direct_55, multiplication_direct_56, multiplication_direct_57, multiplication_direct_58, multiplication_direct_59, multiplication_direct_60, multiplication_direct_61, multiplication_direct_62, multiplication_direct_63, multiplication_direct_64, multiplication_direct_65, multiplication_direct_66, multiplication_direct_67, multiplication_direct_68, multiplication_direct_69,
multiplication_direct_71, multiplication_direct_72, multiplication_direct_73, multiplication_direct_74, multiplication_direct_75, multiplication_direct_76, multiplication_direct_77, multiplication_direct_78, multiplication_direct_79, multiplication_direct_80, multiplication_direct_81, multiplication_direct_82, multiplication_direct_83, multiplication_direct_84, multiplication_direct_85, multiplication_direct_86, multiplication_direct_87, multiplication_direct_88, multiplication_direct_89, multiplication_direct_90, multiplication_direct_91, multiplication_direct_92, multiplication_direct_93, multiplication_direct_94, multiplication_direct_95, multiplication_direct_96, multiplication_direct_97, multiplication_direct_98, multiplication_direct_99, multiplication_direct_100,
multiplication_direct_102, multiplication_direct_103, multiplication_direct_104, multiplication_direct_105, multiplication_direct_106, multiplication_direct_107, multiplication_direct_108, multiplication_direct_109, multiplication_direct_110, multiplication_direct_111, multiplication_direct_112, multiplication_direct_113, multiplication_direct_114, multiplication_direct_115, multiplication_direct_116, multiplication_direct_117, multiplication_direct_118, multiplication_direct_119, multiplication_direct_120, multiplication_direct_121, multiplication_direct_122, multiplication_direct_123, multiplication_direct_124, multiplication_direct_125, multiplication_direct_126, multiplication_direct_127, multiplication_direct_128, multiplication_direct_129, multiplication_direct_130, multiplication_direct_131, multiplication_direct_132, multiplication_direct_133, multiplication_direct_134, multiplication_direct_135, multiplication_direct_136, multiplication_direct_137, multiplication_direct_138, multiplication_direct_139,
-- 0001 square with no reduction
square_direct_0,
square_direct_2, square_direct_3, square_direct_4,
square_direct_6, square_direct_7, square_direct_8, square_direct_9, square_direct_10,
square_direct_12, square_direct_13, square_direct_14, square_direct_15, square_direct_16, square_direct_17, square_direct_18,
square_direct_20, square_direct_21, square_direct_22, square_direct_23, square_direct_24, square_direct_25, square_direct_26, square_direct_27, square_direct_28, square_direct_29,
square_direct_31, square_direct_32, square_direct_33, square_direct_34, square_direct_35, square_direct_36, square_direct_37, square_direct_38, square_direct_39, square_direct_40, square_direct_41, square_direct_42, square_direct_43,
square_direct_45, square_direct_46, square_direct_47, square_direct_48, square_direct_49, square_direct_50, square_direct_51, square_direct_52, square_direct_53, square_direct_54, square_direct_55, square_direct_56, square_direct_57, square_direct_58, square_direct_59, square_direct_60, square_direct_61,
square_direct_63, square_direct_64, square_direct_65, square_direct_66, square_direct_67, square_direct_68, square_direct_69, square_direct_70, square_direct_71, square_direct_72, square_direct_73, square_direct_74, square_direct_75, square_direct_76, square_direct_77, square_direct_78, square_direct_79, square_direct_80, square_direct_81, square_direct_82, square_direct_83,
-- 0010 multiplication with reduction and prime line not equal to 1
multiplication_with_reduction_0, multiplication_with_reduction_1, multiplication_with_reduction_2, multiplication_with_reduction_3,
multiplication_with_reduction_5, multiplication_with_reduction_6, multiplication_with_reduction_7, multiplication_with_reduction_8, multiplication_with_reduction_9, multiplication_with_reduction_10, multiplication_with_reduction_11, multiplication_with_reduction_12, multiplication_with_reduction_13, multiplication_with_reduction_14,
multiplication_with_reduction_16, multiplication_with_reduction_17, multiplication_with_reduction_18, multiplication_with_reduction_19, multiplication_with_reduction_20, multiplication_with_reduction_21, multiplication_with_reduction_22, multiplication_with_reduction_23, multiplication_with_reduction_24, multiplication_with_reduction_25, multiplication_with_reduction_26, multiplication_with_reduction_27, multiplication_with_reduction_28, multiplication_with_reduction_29, multiplication_with_reduction_30, multiplication_with_reduction_31, multiplication_with_reduction_32,
multiplication_with_reduction_34, multiplication_with_reduction_35, multiplication_with_reduction_36, multiplication_with_reduction_37, multiplication_with_reduction_38, multiplication_with_reduction_39, multiplication_with_reduction_40, multiplication_with_reduction_41, multiplication_with_reduction_42, multiplication_with_reduction_43, multiplication_with_reduction_44, multiplication_with_reduction_45, multiplication_with_reduction_46, multiplication_with_reduction_47, multiplication_with_reduction_48, multiplication_with_reduction_49, multiplication_with_reduction_50, multiplication_with_reduction_51, multiplication_with_reduction_52, multiplication_with_reduction_53, multiplication_with_reduction_54, multiplication_with_reduction_55, multiplication_with_reduction_56, multiplication_with_reduction_57, multiplication_with_reduction_58, 
multiplication_with_reduction_60, multiplication_with_reduction_61, multiplication_with_reduction_62, multiplication_with_reduction_63, multiplication_with_reduction_64,multiplication_with_reduction_65, multiplication_with_reduction_66, multiplication_with_reduction_67, multiplication_with_reduction_68, multiplication_with_reduction_69, multiplication_with_reduction_70, multiplication_with_reduction_71, multiplication_with_reduction_72, multiplication_with_reduction_73, multiplication_with_reduction_74,multiplication_with_reduction_75, multiplication_with_reduction_76, multiplication_with_reduction_77, multiplication_with_reduction_78, multiplication_with_reduction_79, multiplication_with_reduction_80, multiplication_with_reduction_81, multiplication_with_reduction_82, multiplication_with_reduction_83, multiplication_with_reduction_84, multiplication_with_reduction_85, multiplication_with_reduction_86, multiplication_with_reduction_87, multiplication_with_reduction_88, multiplication_with_reduction_89, multiplication_with_reduction_90, multiplication_with_reduction_91, multiplication_with_reduction_92, multiplication_with_reduction_93, multiplication_with_reduction_94, multiplication_with_reduction_96, multiplication_with_reduction_97, multiplication_with_reduction_98, multiplication_with_reduction_99, multiplication_with_reduction_100, multiplication_with_reduction_101, multiplication_with_reduction_102, multiplication_with_reduction_103, multiplication_with_reduction_104, multiplication_with_reduction_105, multiplication_with_reduction_106, multiplication_with_reduction_107, multiplication_with_reduction_108, multiplication_with_reduction_109, multiplication_with_reduction_110, multiplication_with_reduction_111, multiplication_with_reduction_112, multiplication_with_reduction_113, multiplication_with_reduction_114, multiplication_with_reduction_115, multiplication_with_reduction_116, multiplication_with_reduction_117, multiplication_with_reduction_118, multiplication_with_reduction_119, multiplication_with_reduction_120, multiplication_with_reduction_121, multiplication_with_reduction_122, multiplication_with_reduction_123, multiplication_with_reduction_124, multiplication_with_reduction_125, multiplication_with_reduction_126, multiplication_with_reduction_127, multiplication_with_reduction_128, multiplication_with_reduction_129, multiplication_with_reduction_130, multiplication_with_reduction_131, multiplication_with_reduction_132, multiplication_with_reduction_133, multiplication_with_reduction_134, multiplication_with_reduction_135, multiplication_with_reduction_136, multiplication_with_reduction_137, multiplication_with_reduction_138, multiplication_with_reduction_139, multiplication_with_reduction_140, multiplication_with_reduction_141, multiplication_with_reduction_142,
multiplication_with_reduction_144, multiplication_with_reduction_145, multiplication_with_reduction_146, multiplication_with_reduction_147, multiplication_with_reduction_148, multiplication_with_reduction_149, multiplication_with_reduction_150, multiplication_with_reduction_151, multiplication_with_reduction_152, multiplication_with_reduction_153, multiplication_with_reduction_154, multiplication_with_reduction_155, multiplication_with_reduction_156, multiplication_with_reduction_157, multiplication_with_reduction_158, multiplication_with_reduction_159, multiplication_with_reduction_160, multiplication_with_reduction_161, multiplication_with_reduction_162, multiplication_with_reduction_163, multiplication_with_reduction_164, multiplication_with_reduction_165, multiplication_with_reduction_166, multiplication_with_reduction_167, multiplication_with_reduction_168, multiplication_with_reduction_169, multiplication_with_reduction_170, multiplication_with_reduction_171, multiplication_with_reduction_172, multiplication_with_reduction_173, multiplication_with_reduction_174, multiplication_with_reduction_175, multiplication_with_reduction_176, multiplication_with_reduction_177, multiplication_with_reduction_178, multiplication_with_reduction_179, multiplication_with_reduction_180, multiplication_with_reduction_181, multiplication_with_reduction_182, multiplication_with_reduction_183, multiplication_with_reduction_184, multiplication_with_reduction_185, multiplication_with_reduction_186, multiplication_with_reduction_187, multiplication_with_reduction_188, multiplication_with_reduction_189, multiplication_with_reduction_190, multiplication_with_reduction_191, multiplication_with_reduction_192, multiplication_with_reduction_193, multiplication_with_reduction_194, multiplication_with_reduction_195, multiplication_with_reduction_196, multiplication_with_reduction_197, multiplication_with_reduction_198, multiplication_with_reduction_199, multiplication_with_reduction_200, multiplication_with_reduction_201, multiplication_with_reduction_202, multiplication_with_reduction_203, multiplication_with_reduction_204,
multiplication_with_reduction_206, multiplication_with_reduction_207, multiplication_with_reduction_208, multiplication_with_reduction_209, multiplication_with_reduction_210, multiplication_with_reduction_211, multiplication_with_reduction_212, multiplication_with_reduction_213, multiplication_with_reduction_214, multiplication_with_reduction_215, multiplication_with_reduction_216, multiplication_with_reduction_217, multiplication_with_reduction_218, multiplication_with_reduction_219, multiplication_with_reduction_220, multiplication_with_reduction_221, multiplication_with_reduction_222, multiplication_with_reduction_223, multiplication_with_reduction_224, multiplication_with_reduction_225, multiplication_with_reduction_226, multiplication_with_reduction_227, multiplication_with_reduction_228, multiplication_with_reduction_229, multiplication_with_reduction_230, multiplication_with_reduction_231, multiplication_with_reduction_232, multiplication_with_reduction_233, multiplication_with_reduction_234, multiplication_with_reduction_235, multiplication_with_reduction_236, multiplication_with_reduction_237, multiplication_with_reduction_238, multiplication_with_reduction_239, multiplication_with_reduction_240, multiplication_with_reduction_241, multiplication_with_reduction_242, multiplication_with_reduction_243, multiplication_with_reduction_244, multiplication_with_reduction_245, multiplication_with_reduction_246, multiplication_with_reduction_247, multiplication_with_reduction_248, multiplication_with_reduction_249, multiplication_with_reduction_250,multiplication_with_reduction_251, multiplication_with_reduction_252, multiplication_with_reduction_253, multiplication_with_reduction_254, multiplication_with_reduction_255, multiplication_with_reduction_256, multiplication_with_reduction_257, multiplication_with_reduction_258, multiplication_with_reduction_259, multiplication_with_reduction_260, multiplication_with_reduction_261, multiplication_with_reduction_262, multiplication_with_reduction_263, multiplication_with_reduction_264, multiplication_with_reduction_265, multiplication_with_reduction_266, multiplication_with_reduction_267, multiplication_with_reduction_268, multiplication_with_reduction_269, multiplication_with_reduction_270, multiplication_with_reduction_271, multiplication_with_reduction_272, multiplication_with_reduction_273, multiplication_with_reduction_274, multiplication_with_reduction_275, multiplication_with_reduction_276, multiplication_with_reduction_277, multiplication_with_reduction_278, multiplication_with_reduction_279, multiplication_with_reduction_280, multiplication_with_reduction_281, multiplication_with_reduction_282,
-- 0010 multiplication with reduction and prime line equal to 1
multiplication_with_reduction_special_prime_0, multiplication_with_reduction_special_prime_1,
multiplication_with_reduction_special_prime_3, multiplication_with_reduction_special_prime_4, multiplication_with_reduction_special_prime_5, multiplication_with_reduction_special_prime_6, multiplication_with_reduction_special_prime_7, multiplication_with_reduction_special_prime_8,
multiplication_with_reduction_special_prime_10, multiplication_with_reduction_special_prime_11, multiplication_with_reduction_special_prime_12, multiplication_with_reduction_special_prime_13, multiplication_with_reduction_special_prime_14, multiplication_with_reduction_special_prime_15, multiplication_with_reduction_special_prime_16, multiplication_with_reduction_special_prime_17, multiplication_with_reduction_special_prime_18, multiplication_with_reduction_special_prime_19, multiplication_with_reduction_special_prime_20,multiplication_with_reduction_special_prime_21, multiplication_with_reduction_special_prime_22, multiplication_with_reduction_special_prime_23,
multiplication_with_reduction_special_prime_25, multiplication_with_reduction_special_prime_26, multiplication_with_reduction_special_prime_27, multiplication_with_reduction_special_prime_28, multiplication_with_reduction_special_prime_29, multiplication_with_reduction_special_prime_30, multiplication_with_reduction_special_prime_31, multiplication_with_reduction_special_prime_32, multiplication_with_reduction_special_prime_33, multiplication_with_reduction_special_prime_34, multiplication_with_reduction_special_prime_35, multiplication_with_reduction_special_prime_36, multiplication_with_reduction_special_prime_37, multiplication_with_reduction_special_prime_38, multiplication_with_reduction_special_prime_39, multiplication_with_reduction_special_prime_40, multiplication_with_reduction_special_prime_41, multiplication_with_reduction_special_prime_42, multiplication_with_reduction_special_prime_43, multiplication_with_reduction_special_prime_44, multiplication_with_reduction_special_prime_45,
multiplication_with_reduction_special_prime_47, multiplication_with_reduction_special_prime_48, multiplication_with_reduction_special_prime_49, multiplication_with_reduction_special_prime_50, multiplication_with_reduction_special_prime_51, multiplication_with_reduction_special_prime_52, multiplication_with_reduction_special_prime_53, multiplication_with_reduction_special_prime_54, multiplication_with_reduction_special_prime_55, multiplication_with_reduction_special_prime_56, multiplication_with_reduction_special_prime_57, multiplication_with_reduction_special_prime_58, multiplication_with_reduction_special_prime_59, multiplication_with_reduction_special_prime_60, multiplication_with_reduction_special_prime_61, multiplication_with_reduction_special_prime_62, multiplication_with_reduction_special_prime_63, multiplication_with_reduction_special_prime_64, multiplication_with_reduction_special_prime_65, multiplication_with_reduction_special_prime_66, multiplication_with_reduction_special_prime_67, multiplication_with_reduction_special_prime_68, multiplication_with_reduction_special_prime_69, multiplication_with_reduction_special_prime_70, multiplication_with_reduction_special_prime_71, multiplication_with_reduction_special_prime_72, multiplication_with_reduction_special_prime_73, multiplication_with_reduction_special_prime_74, multiplication_with_reduction_special_prime_75, multiplication_with_reduction_special_prime_76, multiplication_with_reduction_special_prime_77, multiplication_with_reduction_special_prime_78, multiplication_with_reduction_special_prime_79, multiplication_with_reduction_special_prime_80, multiplication_with_reduction_special_prime_81, multiplication_with_reduction_special_prime_82, multiplication_with_reduction_special_prime_83, multiplication_with_reduction_special_prime_84, multiplication_with_reduction_special_prime_85, multiplication_with_reduction_special_prime_86,
multiplication_with_reduction_special_prime_88, multiplication_with_reduction_special_prime_89, multiplication_with_reduction_special_prime_90, multiplication_with_reduction_special_prime_91, multiplication_with_reduction_special_prime_92, multiplication_with_reduction_special_prime_93, multiplication_with_reduction_special_prime_94, multiplication_with_reduction_special_prime_95, multiplication_with_reduction_special_prime_96, multiplication_with_reduction_special_prime_97, multiplication_with_reduction_special_prime_98, multiplication_with_reduction_special_prime_99, multiplication_with_reduction_special_prime_100, multiplication_with_reduction_special_prime_101, multiplication_with_reduction_special_prime_102, multiplication_with_reduction_special_prime_103, multiplication_with_reduction_special_prime_104, multiplication_with_reduction_special_prime_105, multiplication_with_reduction_special_prime_106, multiplication_with_reduction_special_prime_107, multiplication_with_reduction_special_prime_108, multiplication_with_reduction_special_prime_109, multiplication_with_reduction_special_prime_110, multiplication_with_reduction_special_prime_111, multiplication_with_reduction_special_prime_112, multiplication_with_reduction_special_prime_113, multiplication_with_reduction_special_prime_114, multiplication_with_reduction_special_prime_115, multiplication_with_reduction_special_prime_116, multiplication_with_reduction_special_prime_117, multiplication_with_reduction_special_prime_118, multiplication_with_reduction_special_prime_119, multiplication_with_reduction_special_prime_120, multiplication_with_reduction_special_prime_121, multiplication_with_reduction_special_prime_122, multiplication_with_reduction_special_prime_123, multiplication_with_reduction_special_prime_124, multiplication_with_reduction_special_prime_125, multiplication_with_reduction_special_prime_126, multiplication_with_reduction_special_prime_127, multiplication_with_reduction_special_prime_128,
multiplication_with_reduction_special_prime_130, multiplication_with_reduction_special_prime_131, multiplication_with_reduction_special_prime_132, multiplication_with_reduction_special_prime_133, multiplication_with_reduction_special_prime_134, multiplication_with_reduction_special_prime_135, multiplication_with_reduction_special_prime_136, multiplication_with_reduction_special_prime_137, multiplication_with_reduction_special_prime_138, multiplication_with_reduction_special_prime_139, multiplication_with_reduction_special_prime_140, multiplication_with_reduction_special_prime_141, multiplication_with_reduction_special_prime_142, multiplication_with_reduction_special_prime_143, multiplication_with_reduction_special_prime_144, multiplication_with_reduction_special_prime_145, multiplication_with_reduction_special_prime_146, multiplication_with_reduction_special_prime_147, multiplication_with_reduction_special_prime_148, multiplication_with_reduction_special_prime_149, multiplication_with_reduction_special_prime_150, multiplication_with_reduction_special_prime_151, multiplication_with_reduction_special_prime_152, multiplication_with_reduction_special_prime_153, multiplication_with_reduction_special_prime_154, multiplication_with_reduction_special_prime_155, multiplication_with_reduction_special_prime_156, multiplication_with_reduction_special_prime_157, multiplication_with_reduction_special_prime_158, multiplication_with_reduction_special_prime_159, multiplication_with_reduction_special_prime_160, multiplication_with_reduction_special_prime_161, multiplication_with_reduction_special_prime_162, multiplication_with_reduction_special_prime_163, multiplication_with_reduction_special_prime_164, multiplication_with_reduction_special_prime_165, multiplication_with_reduction_special_prime_166, multiplication_with_reduction_special_prime_167, multiplication_with_reduction_special_prime_168, multiplication_with_reduction_special_prime_169, multiplication_with_reduction_special_prime_170, multiplication_with_reduction_special_prime_171, multiplication_with_reduction_special_prime_172, multiplication_with_reduction_special_prime_173, multiplication_with_reduction_special_prime_174, multiplication_with_reduction_special_prime_175, multiplication_with_reduction_special_prime_176, multiplication_with_reduction_special_prime_177, multiplication_with_reduction_special_prime_178, multiplication_with_reduction_special_prime_179, multiplication_with_reduction_special_prime_180, multiplication_with_reduction_special_prime_181, multiplication_with_reduction_special_prime_182, multiplication_with_reduction_special_prime_183, multiplication_with_reduction_special_prime_184, multiplication_with_reduction_special_prime_185, multiplication_with_reduction_special_prime_186, multiplication_with_reduction_special_prime_187, multiplication_with_reduction_special_prime_188, multiplication_with_reduction_special_prime_189, multiplication_with_reduction_special_prime_190, multiplication_with_reduction_special_prime_191, multiplication_with_reduction_special_prime_192, multiplication_with_reduction_special_prime_193, multiplication_with_reduction_special_prime_194, multiplication_with_reduction_special_prime_195, multiplication_with_reduction_special_prime_196, multiplication_with_reduction_special_prime_197, multiplication_with_reduction_special_prime_198, multiplication_with_reduction_special_prime_199, multiplication_with_reduction_special_prime_200, multiplication_with_reduction_special_prime_201, multiplication_with_reduction_special_prime_202, multiplication_with_reduction_special_prime_203, multiplication_with_reduction_special_prime_204, multiplication_with_reduction_special_prime_205, multiplication_with_reduction_special_prime_206,
multiplication_with_reduction_special_prime_208, multiplication_with_reduction_special_prime_209, multiplication_with_reduction_special_prime_210, multiplication_with_reduction_special_prime_211, multiplication_with_reduction_special_prime_212, multiplication_with_reduction_special_prime_213, multiplication_with_reduction_special_prime_214, multiplication_with_reduction_special_prime_215, multiplication_with_reduction_special_prime_216, multiplication_with_reduction_special_prime_217, multiplication_with_reduction_special_prime_218, multiplication_with_reduction_special_prime_219, multiplication_with_reduction_special_prime_220, multiplication_with_reduction_special_prime_221, multiplication_with_reduction_special_prime_222, multiplication_with_reduction_special_prime_223, multiplication_with_reduction_special_prime_224, multiplication_with_reduction_special_prime_225, multiplication_with_reduction_special_prime_226, multiplication_with_reduction_special_prime_227, multiplication_with_reduction_special_prime_228, multiplication_with_reduction_special_prime_229, multiplication_with_reduction_special_prime_230, multiplication_with_reduction_special_prime_231, multiplication_with_reduction_special_prime_232, multiplication_with_reduction_special_prime_233, multiplication_with_reduction_special_prime_234, multiplication_with_reduction_special_prime_235, multiplication_with_reduction_special_prime_236, multiplication_with_reduction_special_prime_237, multiplication_with_reduction_special_prime_238, multiplication_with_reduction_special_prime_239, multiplication_with_reduction_special_prime_240, multiplication_with_reduction_special_prime_241, multiplication_with_reduction_special_prime_242, multiplication_with_reduction_special_prime_243, multiplication_with_reduction_special_prime_244, multiplication_with_reduction_special_prime_245, multiplication_with_reduction_special_prime_246, multiplication_with_reduction_special_prime_247, multiplication_with_reduction_special_prime_248, multiplication_with_reduction_special_prime_249, multiplication_with_reduction_special_prime_250, multiplication_with_reduction_special_prime_251, multiplication_with_reduction_special_prime_252, multiplication_with_reduction_special_prime_253, multiplication_with_reduction_special_prime_254, multiplication_with_reduction_special_prime_255, multiplication_with_reduction_special_prime_256, multiplication_with_reduction_special_prime_257, multiplication_with_reduction_special_prime_258, multiplication_with_reduction_special_prime_259, multiplication_with_reduction_special_prime_260, multiplication_with_reduction_special_prime_261, multiplication_with_reduction_special_prime_262, multiplication_with_reduction_special_prime_263, multiplication_with_reduction_special_prime_264, multiplication_with_reduction_special_prime_265, multiplication_with_reduction_special_prime_266, multiplication_with_reduction_special_prime_267, multiplication_with_reduction_special_prime_268, multiplication_with_reduction_special_prime_269, multiplication_with_reduction_special_prime_270, multiplication_with_reduction_special_prime_271, multiplication_with_reduction_special_prime_272, multiplication_with_reduction_special_prime_273, multiplication_with_reduction_special_prime_274, multiplication_with_reduction_special_prime_275,
-- 0011 square with reduction and prime line not equal to 1
square_with_reduction_0, square_with_reduction_1, square_with_reduction_2, square_with_reduction_3,
square_with_reduction_5, square_with_reduction_6, square_with_reduction_7, square_with_reduction_8, square_with_reduction_9, square_with_reduction_10, square_with_reduction_11, square_with_reduction_12, square_with_reduction_13,
square_with_reduction_15, square_with_reduction_16, square_with_reduction_17, square_with_reduction_18, square_with_reduction_19, square_with_reduction_20, square_with_reduction_21, square_with_reduction_22, square_with_reduction_23, square_with_reduction_24, square_with_reduction_25, square_with_reduction_26, square_with_reduction_27, square_with_reduction_28, 
square_with_reduction_30, square_with_reduction_31, square_with_reduction_32, square_with_reduction_33, square_with_reduction_34, square_with_reduction_35, square_with_reduction_36, square_with_reduction_37, square_with_reduction_38, square_with_reduction_39, square_with_reduction_40, square_with_reduction_41, square_with_reduction_42, square_with_reduction_43, square_with_reduction_44, square_with_reduction_45, square_with_reduction_46, square_with_reduction_47, square_with_reduction_48, square_with_reduction_49,
square_with_reduction_51, square_with_reduction_52, square_with_reduction_53, square_with_reduction_54, square_with_reduction_55, square_with_reduction_56, square_with_reduction_57, square_with_reduction_58, square_with_reduction_59, square_with_reduction_60, square_with_reduction_61, square_with_reduction_62, square_with_reduction_63, square_with_reduction_64, square_with_reduction_65, square_with_reduction_66, square_with_reduction_67, square_with_reduction_68, square_with_reduction_69, square_with_reduction_70, square_with_reduction_71, square_with_reduction_72, square_with_reduction_73, square_with_reduction_74, square_with_reduction_75, square_with_reduction_76, square_with_reduction_77, square_with_reduction_78,
square_with_reduction_80, square_with_reduction_81, square_with_reduction_82, square_with_reduction_83, square_with_reduction_84, square_with_reduction_85, square_with_reduction_86, square_with_reduction_87, square_with_reduction_88, square_with_reduction_89, square_with_reduction_90, square_with_reduction_91, square_with_reduction_92, square_with_reduction_93, square_with_reduction_94, square_with_reduction_95, square_with_reduction_96, square_with_reduction_97, square_with_reduction_98, square_with_reduction_99, square_with_reduction_100, square_with_reduction_101, square_with_reduction_102, square_with_reduction_103, square_with_reduction_104, square_with_reduction_105, square_with_reduction_106, square_with_reduction_107, square_with_reduction_108, square_with_reduction_109, square_with_reduction_110, square_with_reduction_111, square_with_reduction_112, square_with_reduction_113, square_with_reduction_114, square_with_reduction_115, square_with_reduction_116,
square_with_reduction_118, square_with_reduction_119, square_with_reduction_120, square_with_reduction_121, square_with_reduction_122, square_with_reduction_123, square_with_reduction_124, square_with_reduction_125, square_with_reduction_126, square_with_reduction_127, square_with_reduction_128, square_with_reduction_129, square_with_reduction_130, square_with_reduction_131, square_with_reduction_132, square_with_reduction_133, square_with_reduction_134, square_with_reduction_135, square_with_reduction_136, square_with_reduction_137, square_with_reduction_138, square_with_reduction_139, square_with_reduction_140, square_with_reduction_141, square_with_reduction_142, square_with_reduction_143, square_with_reduction_144, square_with_reduction_145, square_with_reduction_146, square_with_reduction_147, square_with_reduction_148, square_with_reduction_149, square_with_reduction_150, square_with_reduction_151, square_with_reduction_152, square_with_reduction_153, square_with_reduction_154, square_with_reduction_155, square_with_reduction_156, square_with_reduction_157, square_with_reduction_158, square_with_reduction_159, square_with_reduction_160, square_with_reduction_161, square_with_reduction_162, square_with_reduction_163, square_with_reduction_164, square_with_reduction_165,
square_with_reduction_167, square_with_reduction_168, square_with_reduction_169, square_with_reduction_170, square_with_reduction_171, square_with_reduction_172, square_with_reduction_173, square_with_reduction_174, square_with_reduction_175, square_with_reduction_176, square_with_reduction_177, square_with_reduction_178, square_with_reduction_179, square_with_reduction_180, square_with_reduction_181, square_with_reduction_182, square_with_reduction_183, square_with_reduction_184, square_with_reduction_185, square_with_reduction_186, square_with_reduction_187, square_with_reduction_188, square_with_reduction_189, square_with_reduction_190, square_with_reduction_191, square_with_reduction_192, square_with_reduction_193, square_with_reduction_194, square_with_reduction_195, square_with_reduction_196, square_with_reduction_197, square_with_reduction_198, square_with_reduction_199, square_with_reduction_200, square_with_reduction_201, square_with_reduction_202, square_with_reduction_203, square_with_reduction_204, square_with_reduction_205, square_with_reduction_206, square_with_reduction_207, square_with_reduction_208, square_with_reduction_209, square_with_reduction_210, square_with_reduction_211, square_with_reduction_212, square_with_reduction_213, square_with_reduction_214, square_with_reduction_215, square_with_reduction_216, square_with_reduction_217, square_with_reduction_218, square_with_reduction_219, square_with_reduction_220, square_with_reduction_221, square_with_reduction_222, square_with_reduction_223, square_with_reduction_224, square_with_reduction_225, square_with_reduction_226,
-- 0011 square with reduction and prime line equal to 1
square_with_reduction_special_prime_0, square_with_reduction_special_prime_1,
square_with_reduction_special_prime_3, square_with_reduction_special_prime_4, square_with_reduction_special_prime_5, square_with_reduction_special_prime_6, square_with_reduction_special_prime_7,
square_with_reduction_special_prime_9, square_with_reduction_special_prime_10, square_with_reduction_special_prime_11, square_with_reduction_special_prime_12, square_with_reduction_special_prime_13, square_with_reduction_special_prime_14, square_with_reduction_special_prime_15, square_with_reduction_special_prime_16, square_with_reduction_special_prime_17, square_with_reduction_special_prime_18,
square_with_reduction_special_prime_20, square_with_reduction_special_prime_21, square_with_reduction_special_prime_22, square_with_reduction_special_prime_23, square_with_reduction_special_prime_24, square_with_reduction_special_prime_25, square_with_reduction_special_prime_26, square_with_reduction_special_prime_27, square_with_reduction_special_prime_28, square_with_reduction_special_prime_29, square_with_reduction_special_prime_30, square_with_reduction_special_prime_31, square_with_reduction_special_prime_32, square_with_reduction_special_prime_33, square_with_reduction_special_prime_34, square_with_reduction_special_prime_35, 
square_with_reduction_special_prime_37, square_with_reduction_special_prime_38, square_with_reduction_special_prime_39, square_with_reduction_special_prime_40, square_with_reduction_special_prime_41, square_with_reduction_special_prime_42, square_with_reduction_special_prime_43, square_with_reduction_special_prime_44, square_with_reduction_special_prime_45, square_with_reduction_special_prime_46, square_with_reduction_special_prime_47, square_with_reduction_special_prime_48, square_with_reduction_special_prime_49, square_with_reduction_special_prime_50, square_with_reduction_special_prime_51, square_with_reduction_special_prime_52, square_with_reduction_special_prime_53, square_with_reduction_special_prime_54, square_with_reduction_special_prime_55, square_with_reduction_special_prime_56, square_with_reduction_special_prime_57, square_with_reduction_special_prime_58, square_with_reduction_special_prime_59, square_with_reduction_special_prime_60, square_with_reduction_special_prime_61, square_with_reduction_special_prime_62, square_with_reduction_special_prime_63, square_with_reduction_special_prime_64, square_with_reduction_special_prime_65, square_with_reduction_special_prime_66,
square_with_reduction_special_prime_68, square_with_reduction_special_prime_69, square_with_reduction_special_prime_70, square_with_reduction_special_prime_71, square_with_reduction_special_prime_72, square_with_reduction_special_prime_73, square_with_reduction_special_prime_74, square_with_reduction_special_prime_75, square_with_reduction_special_prime_76, square_with_reduction_special_prime_77, square_with_reduction_special_prime_78, square_with_reduction_special_prime_79, square_with_reduction_special_prime_80, square_with_reduction_special_prime_81, square_with_reduction_special_prime_82, square_with_reduction_special_prime_83, square_with_reduction_special_prime_84, square_with_reduction_special_prime_85, square_with_reduction_special_prime_86, square_with_reduction_special_prime_87, square_with_reduction_special_prime_88, square_with_reduction_special_prime_89, square_with_reduction_special_prime_90, square_with_reduction_special_prime_91, square_with_reduction_special_prime_92, square_with_reduction_special_prime_93, square_with_reduction_special_prime_94, square_with_reduction_special_prime_95, square_with_reduction_special_prime_96, square_with_reduction_special_prime_97, square_with_reduction_special_prime_98,
square_with_reduction_special_prime_100, square_with_reduction_special_prime_101, square_with_reduction_special_prime_102, square_with_reduction_special_prime_103, square_with_reduction_special_prime_104, square_with_reduction_special_prime_105, square_with_reduction_special_prime_106, square_with_reduction_special_prime_107, square_with_reduction_special_prime_108, square_with_reduction_special_prime_109, square_with_reduction_special_prime_110, square_with_reduction_special_prime_111, square_with_reduction_special_prime_112, square_with_reduction_special_prime_113, square_with_reduction_special_prime_114, square_with_reduction_special_prime_115, square_with_reduction_special_prime_116, square_with_reduction_special_prime_117, square_with_reduction_special_prime_118, square_with_reduction_special_prime_119, square_with_reduction_special_prime_120, square_with_reduction_special_prime_121, square_with_reduction_special_prime_122, square_with_reduction_special_prime_123, square_with_reduction_special_prime_124, square_with_reduction_special_prime_125, square_with_reduction_special_prime_126, square_with_reduction_special_prime_127, square_with_reduction_special_prime_128, square_with_reduction_special_prime_129, square_with_reduction_special_prime_130, square_with_reduction_special_prime_131, square_with_reduction_special_prime_132, square_with_reduction_special_prime_133, square_with_reduction_special_prime_134, square_with_reduction_special_prime_135, square_with_reduction_special_prime_136, square_with_reduction_special_prime_137, square_with_reduction_special_prime_138, square_with_reduction_special_prime_139, square_with_reduction_special_prime_140, square_with_reduction_special_prime_141, square_with_reduction_special_prime_142, square_with_reduction_special_prime_143, square_with_reduction_special_prime_144, square_with_reduction_special_prime_145, square_with_reduction_special_prime_146, square_with_reduction_special_prime_147, square_with_reduction_special_prime_148, square_with_reduction_special_prime_149, square_with_reduction_special_prime_150, square_with_reduction_special_prime_151, square_with_reduction_special_prime_152, square_with_reduction_special_prime_153, square_with_reduction_special_prime_154, square_with_reduction_special_prime_155,
square_with_reduction_special_prime_157, square_with_reduction_special_prime_158, square_with_reduction_special_prime_159, square_with_reduction_special_prime_160, square_with_reduction_special_prime_161, square_with_reduction_special_prime_162, square_with_reduction_special_prime_163, square_with_reduction_special_prime_164, square_with_reduction_special_prime_165, square_with_reduction_special_prime_166, square_with_reduction_special_prime_167, square_with_reduction_special_prime_168, square_with_reduction_special_prime_169, square_with_reduction_special_prime_170, square_with_reduction_special_prime_171, square_with_reduction_special_prime_172, square_with_reduction_special_prime_173, square_with_reduction_special_prime_174, square_with_reduction_special_prime_175, square_with_reduction_special_prime_176, square_with_reduction_special_prime_177, square_with_reduction_special_prime_178, square_with_reduction_special_prime_179, square_with_reduction_special_prime_180, square_with_reduction_special_prime_181, square_with_reduction_special_prime_182, square_with_reduction_special_prime_183, square_with_reduction_special_prime_184, square_with_reduction_special_prime_185, square_with_reduction_special_prime_186, square_with_reduction_special_prime_187, square_with_reduction_special_prime_188, square_with_reduction_special_prime_189, square_with_reduction_special_prime_190, square_with_reduction_special_prime_191, square_with_reduction_special_prime_192, square_with_reduction_special_prime_193, square_with_reduction_special_prime_194, square_with_reduction_special_prime_195, square_with_reduction_special_prime_196, square_with_reduction_special_prime_197, square_with_reduction_special_prime_198, square_with_reduction_special_prime_199, square_with_reduction_special_prime_200, square_with_reduction_special_prime_201, square_with_reduction_special_prime_202, square_with_reduction_special_prime_203, square_with_reduction_special_prime_204, square_with_reduction_special_prime_205, square_with_reduction_special_prime_206, square_with_reduction_special_prime_207,
-- 0100 addition with no reduction
addition_subtraction_direct_0, addition_subtraction_direct_2, addition_subtraction_direct_3, addition_subtraction_direct_5, addition_subtraction_direct_6, addition_subtraction_direct_8, addition_subtraction_direct_9, addition_subtraction_direct_11, addition_subtraction_direct_12, addition_subtraction_direct_14, addition_subtraction_direct_15, addition_subtraction_direct_17, addition_subtraction_direct_18, addition_subtraction_direct_20, addition_subtraction_direct_21,
-- 0101 iterative modular reduction
iterative_modular_reduction_0, iterative_modular_reduction_1, iterative_modular_reduction_2, iterative_modular_reduction_3,
iterative_modular_reduction_5, iterative_modular_reduction_6, iterative_modular_reduction_7, iterative_modular_reduction_8, iterative_modular_reduction_9, iterative_modular_reduction_10, iterative_modular_reduction_11,
iterative_modular_reduction_13, iterative_modular_reduction_14, iterative_modular_reduction_15, iterative_modular_reduction_16, iterative_modular_reduction_17, iterative_modular_reduction_18, iterative_modular_reduction_19, iterative_modular_reduction_20, iterative_modular_reduction_21, iterative_modular_reduction_22,
iterative_modular_reduction_24, iterative_modular_reduction_25, iterative_modular_reduction_26, iterative_modular_reduction_27, iterative_modular_reduction_28, iterative_modular_reduction_29, iterative_modular_reduction_30, iterative_modular_reduction_31, iterative_modular_reduction_32, iterative_modular_reduction_33, iterative_modular_reduction_34, iterative_modular_reduction_35, iterative_modular_reduction_36,
iterative_modular_reduction_38, iterative_modular_reduction_39, iterative_modular_reduction_40, iterative_modular_reduction_41, iterative_modular_reduction_42, iterative_modular_reduction_43, iterative_modular_reduction_44, iterative_modular_reduction_45, iterative_modular_reduction_46, iterative_modular_reduction_47, iterative_modular_reduction_48, iterative_modular_reduction_49, iterative_modular_reduction_50, iterative_modular_reduction_51, iterative_modular_reduction_52, iterative_modular_reduction_53,
iterative_modular_reduction_55, iterative_modular_reduction_56, iterative_modular_reduction_57, iterative_modular_reduction_58, iterative_modular_reduction_59, iterative_modular_reduction_60, iterative_modular_reduction_61, iterative_modular_reduction_62, iterative_modular_reduction_63, iterative_modular_reduction_64, iterative_modular_reduction_65, iterative_modular_reduction_66, iterative_modular_reduction_67, iterative_modular_reduction_68, iterative_modular_reduction_69, iterative_modular_reduction_70, iterative_modular_reduction_71, iterative_modular_reduction_72, iterative_modular_reduction_73,
iterative_modular_reduction_75, iterative_modular_reduction_76, iterative_modular_reduction_77, iterative_modular_reduction_78, iterative_modular_reduction_79, iterative_modular_reduction_80, iterative_modular_reduction_81, iterative_modular_reduction_82, iterative_modular_reduction_83, iterative_modular_reduction_84, iterative_modular_reduction_85, iterative_modular_reduction_86, iterative_modular_reduction_87, iterative_modular_reduction_88, iterative_modular_reduction_89, iterative_modular_reduction_90, iterative_modular_reduction_91, iterative_modular_reduction_92, iterative_modular_reduction_93, iterative_modular_reduction_94, iterative_modular_reduction_95, iterative_modular_reduction_96,
iterative_modular_reduction_98, iterative_modular_reduction_99, iterative_modular_reduction_100, iterative_modular_reduction_101, iterative_modular_reduction_102, iterative_modular_reduction_103, iterative_modular_reduction_104, iterative_modular_reduction_105, iterative_modular_reduction_106, iterative_modular_reduction_107, iterative_modular_reduction_108, iterative_modular_reduction_109, iterative_modular_reduction_110, iterative_modular_reduction_111, iterative_modular_reduction_112, iterative_modular_reduction_113, iterative_modular_reduction_114, iterative_modular_reduction_115, iterative_modular_reduction_116, iterative_modular_reduction_117, iterative_modular_reduction_118, iterative_modular_reduction_119, iterative_modular_reduction_120, iterative_modular_reduction_121, iterative_modular_reduction_122,
-- NOP
nop_4_stages, nop_8_stages
); 

signal actual_state, next_state : state;

signal next_sm_rotation_size : std_logic_vector(1 downto 0);
signal next_sm_circular_shift_enable : std_logic;
signal next_sel_address_a : std_logic;
signal next_sel_address_b_prime : std_logic_vector(1 downto 0);
signal next_sm_specific_mac_address_a : std_logic_vector(2 downto 0);
signal next_sm_specific_mac_address_b : std_logic_vector(2 downto 0);
signal next_sm_specific_mac_address_o : std_logic_vector(2 downto 0);
signal next_sm_specific_mac_next_address_o : std_logic_vector(2 downto 0);
signal next_mac_enable_signed_a : std_logic;
signal next_mac_enable_signed_b : std_logic;
signal next_mac_sel_load_reg_a : std_logic_vector(1 downto 0);
signal next_mac_clear_reg_b : std_logic;
signal next_mac_clear_reg_acc : std_logic;
signal next_mac_sel_shift_reg_o : std_logic;
signal next_mac_enable_update_reg_s : std_logic;
signal next_mac_sel_reg_s_reg_o_sign : std_logic;
signal next_mac_reg_s_reg_o_positive : std_logic;
signal next_sm_sign_a_mode : std_logic;
signal next_sm_mac_operation_mode : std_logic_vector(1 downto 0);
signal next_mac_enable_reg_s_mask : std_logic;
signal next_mac_subtraction_reg_a_b : std_logic;
signal next_mac_sel_multiply_two_a_b : std_logic;
signal next_mac_sel_reg_y_output : std_logic;
signal next_sm_mac_write_enable_output : std_logic;
signal next_mac_memory_double_mode : std_logic;
signal next_mac_memory_only_write_mode : std_logic;
signal next_base_address_generator_o_increment_previous_address : std_logic;
signal next_sm_free_flag : std_logic;

begin

registers_state : process(clk, rstn)
begin
    if(rstn = '0') then
        actual_state <= reset;
    elsif(rising_edge(clk)) then
        actual_state <= next_state;
    end if;
end process;

registers_state_output : process(clk)
begin
    if(rising_edge(clk)) then
        if(rstn = '0') then
            sm_free_flag <= '0';
            sm_rotation_size <= "11";
            sm_circular_shift_enable <= '0';
            sel_address_a <= '0';
            sel_address_b_prime <= "00";
            sm_specific_mac_address_a <= "000";
            sm_specific_mac_address_b <= "000";
            sm_specific_mac_address_o <= "000";
            sm_specific_mac_next_address_o <= "001";
            mac_enable_signed_a <= '0';
            mac_enable_signed_b <= '0';
            mac_sel_load_reg_a <= "11";
            mac_clear_reg_b <= '1';
            mac_clear_reg_acc <= '1';
            mac_sel_shift_reg_o <= '0';
            mac_enable_update_reg_s <= '0';
            mac_sel_reg_s_reg_o_sign <= '0';
            mac_reg_s_reg_o_positive <= '0';
            sm_sign_a_mode <= '0';
            sm_mac_operation_mode <= "10";
            mac_enable_reg_s_mask <= '0';
            mac_subtraction_reg_a_b <= '0';
            mac_sel_multiply_two_a_b <= '0';
            mac_sel_reg_y_output <= '0';
            base_address_generator_o_increment_previous_address <= '0';
            sm_mac_write_enable_output <= '0';
            mac_memory_double_mode <= '0';
            mac_memory_only_write_mode <= '0';
        else
            sm_free_flag <= next_sm_free_flag;
            sm_rotation_size <= next_sm_rotation_size;
            sm_circular_shift_enable <= next_sm_circular_shift_enable;
            sel_address_a <= next_sel_address_a;
            sel_address_b_prime <= next_sel_address_b_prime;
            sm_specific_mac_address_a <= next_sm_specific_mac_address_a;
            sm_specific_mac_address_b <= next_sm_specific_mac_address_b;
            sm_specific_mac_address_o <= next_sm_specific_mac_address_o;
            sm_specific_mac_next_address_o <= next_sm_specific_mac_next_address_o;
            mac_enable_signed_a <= next_mac_enable_signed_a;
            mac_enable_signed_b <= next_mac_enable_signed_b;
            mac_sel_load_reg_a <= next_mac_sel_load_reg_a;
            mac_clear_reg_b <= next_mac_clear_reg_b;
            mac_clear_reg_acc <= next_mac_clear_reg_acc;
            mac_sel_shift_reg_o <= next_mac_sel_shift_reg_o;
            mac_enable_update_reg_s <= next_mac_enable_update_reg_s;
            mac_sel_reg_s_reg_o_sign <= next_mac_sel_reg_s_reg_o_sign;
            mac_reg_s_reg_o_positive <= next_mac_reg_s_reg_o_positive;
            sm_sign_a_mode <= next_sm_sign_a_mode;
            sm_mac_operation_mode <= next_sm_mac_operation_mode;
            mac_enable_reg_s_mask <= next_mac_enable_reg_s_mask;
            mac_subtraction_reg_a_b <= next_mac_subtraction_reg_a_b;
            mac_sel_multiply_two_a_b <= next_mac_sel_multiply_two_a_b;
            mac_sel_reg_y_output <= next_mac_sel_reg_y_output;
            base_address_generator_o_increment_previous_address <= next_base_address_generator_o_increment_previous_address;
            sm_mac_write_enable_output <= next_sm_mac_write_enable_output;
            mac_memory_double_mode <= next_mac_memory_double_mode;
            mac_memory_only_write_mode <= next_mac_memory_only_write_mode;
        end if;
    end if;
end process;

update_output : process(actual_state, instruction_values_valid, instruction_type, operands_size, prime_line_equal_one)
begin
    case (actual_state) is
        when reset =>
            next_sm_free_flag <= '1';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '0';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "11";
            next_mac_clear_reg_b <= '1';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when decode_instruction =>
            next_sm_free_flag <= '1';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '0';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "11";
            next_mac_clear_reg_b <= '1';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
            if(instruction_values_valid = '1') then
                next_sm_free_flag <= '0';
                if(instruction_type = "0000") then
                    if(operands_size = "000") then
                        -- multiplication_direct_0;
                        -- -- In case of size 1
                        -- reg_a = a0_X; reg_b = b0_X; reg_acc = 0; o0_X = reg_o; o1_X = reg_o >> 272; Enable sign a,b; operation : a*b + acc;
                        next_sm_free_flag <= '0';
                        next_sm_rotation_size <= "11";
                        next_sm_circular_shift_enable <= '1';
                        next_sel_address_a <= '0';
                        next_sel_address_b_prime <= "00";
                        next_sm_specific_mac_address_a <= "000";
                        next_sm_specific_mac_address_b <= "000";
                        next_sm_specific_mac_address_o <= "000";
                        next_sm_specific_mac_next_address_o <= "001";
                        next_mac_enable_signed_a <= '1';
                        next_mac_enable_signed_b <= '1';
                        next_mac_sel_load_reg_a <= "00";
                        next_mac_clear_reg_b <= '0';
                        next_mac_clear_reg_acc <= '1';
                        next_mac_sel_shift_reg_o <= '0';
                        next_mac_enable_update_reg_s <= '0';
                        next_mac_sel_reg_s_reg_o_sign <= '0';
                        next_mac_reg_s_reg_o_positive <= '0';
                        next_sm_sign_a_mode <= '0';
                        next_sm_mac_operation_mode <= "10";
                        next_mac_enable_reg_s_mask <= '0';
                        next_mac_subtraction_reg_a_b <= '0';
                        next_mac_sel_multiply_two_a_b <= '0';
                        next_mac_sel_reg_y_output <= '0';
                        next_sm_mac_write_enable_output <= '1';
                        next_mac_memory_double_mode <= '1';
                        next_mac_memory_only_write_mode <= '1';
                        next_base_address_generator_o_increment_previous_address <= '0';
                    else
                        -- multiplication_direct_2;
                        -- -- Other cases
                        -- reg_a = a0_X; reg_b = b0_X; reg_acc = 0; o0_X = reg_o; operation : a*b + acc; o0_X = reg_o;
                        next_sm_free_flag <= '0';
                        next_sm_rotation_size <= "11";
                        next_sm_circular_shift_enable <= '1';
                        next_sel_address_a <= '0';
                        next_sel_address_b_prime <= "00";
                        next_sm_specific_mac_address_a <= "000";
                        next_sm_specific_mac_address_b <= "000";
                        next_sm_specific_mac_address_o <= "000";
                        next_sm_specific_mac_next_address_o <= "001";
                        next_mac_enable_signed_a <= '0';
                        next_mac_enable_signed_b <= '0';
                        next_mac_sel_load_reg_a <= "00";
                        next_mac_clear_reg_b <= '0';
                        next_mac_clear_reg_acc <= '1';
                        next_mac_sel_shift_reg_o <= '0';
                        next_mac_enable_update_reg_s <= '0';
                        next_mac_sel_reg_s_reg_o_sign <= '0';
                        next_mac_reg_s_reg_o_positive <= '0';
                        next_sm_sign_a_mode <= '0';
                        next_sm_mac_operation_mode <= "10";
                        next_mac_enable_reg_s_mask <= '0';
                        next_mac_subtraction_reg_a_b <= '0';
                        next_mac_sel_multiply_two_a_b <= '0';
                        next_mac_sel_reg_y_output <= '0';
                        next_sm_mac_write_enable_output <= '1';
                        next_mac_memory_double_mode <= '0';
                        next_mac_memory_only_write_mode <= '0';
                        next_base_address_generator_o_increment_previous_address <= '0';
                    end if;
                elsif(instruction_type = "0001") then
                    if(operands_size = "000") then
                        -- square_direct_0;
                        -- -- In case of size 1
                        -- reg_a = a0_X; reg_b = a0_X; reg_acc = 0; o0_X = reg_o; o1_X = reg_o >> 272; Enable sign a,b; operation : a*b + acc;
                        next_sm_free_flag <= '0';
                        next_sm_rotation_size <= "11";
                        next_sm_circular_shift_enable <= '1';
                        next_sel_address_a <= '0';
                        next_sel_address_b_prime <= "00";
                        next_sm_specific_mac_address_a <= "000";
                        next_sm_specific_mac_address_b <= "000";
                        next_sm_specific_mac_address_o <= "000";
                        next_sm_specific_mac_next_address_o <= "001";
                        next_mac_enable_signed_a <= '1';
                        next_mac_enable_signed_b <= '1';
                        next_mac_sel_load_reg_a <= "00";
                        next_mac_clear_reg_b <= '0';
                        next_mac_clear_reg_acc <= '1';
                        next_mac_sel_shift_reg_o <= '0';
                        next_mac_enable_update_reg_s <= '0';
                        next_mac_sel_reg_s_reg_o_sign <= '0';
                        next_mac_reg_s_reg_o_positive <= '0';
                        next_sm_sign_a_mode <= '0';
                        next_sm_mac_operation_mode <= "10";
                        next_mac_enable_reg_s_mask <= '0';
                        next_mac_subtraction_reg_a_b <= '0';
                        next_mac_sel_multiply_two_a_b <= '0';
                        next_mac_sel_reg_y_output <= '0';
                        next_sm_mac_write_enable_output <= '1';
                        next_mac_memory_double_mode <= '1';
                        next_mac_memory_only_write_mode <= '1';
                        next_base_address_generator_o_increment_previous_address <= '0';
                    else
                        -- square_direct_2;
                        -- -- In case of sizes 2, 3, 4, 5, 6, 7, 8
                        -- reg_a = a0_X; reg_b = a0_X; reg_acc = 0; o0_X = reg_o; operation : a*b + acc;
                        next_sm_free_flag <= '0';
                        next_sm_rotation_size <= "11";
                        next_sm_circular_shift_enable <= '1';
                        next_sel_address_a <= '0';
                        next_sel_address_b_prime <= "00";
                        next_sm_specific_mac_address_a <= "000";
                        next_sm_specific_mac_address_b <= "000";
                        next_sm_specific_mac_address_o <= "000";
                        next_sm_specific_mac_next_address_o <= "001";
                        next_mac_enable_signed_a <= '0';
                        next_mac_enable_signed_b <= '0';
                        next_mac_sel_load_reg_a <= "00";
                        next_mac_clear_reg_b <= '0';
                        next_mac_clear_reg_acc <= '1';
                        next_mac_sel_shift_reg_o <= '0';
                        next_mac_enable_update_reg_s <= '0';
                        next_mac_sel_reg_s_reg_o_sign <= '0';
                        next_mac_reg_s_reg_o_positive <= '0';
                        next_sm_sign_a_mode <= '0';
                        next_sm_mac_operation_mode <= "10";
                        next_mac_enable_reg_s_mask <= '0';
                        next_mac_subtraction_reg_a_b <= '0';
                        next_mac_sel_multiply_two_a_b <= '0';
                        next_mac_sel_reg_y_output <= '0';
                        next_sm_mac_write_enable_output <= '1';
                        next_mac_memory_double_mode <= '0';
                        next_mac_memory_only_write_mode <= '0';
                        next_base_address_generator_o_increment_previous_address <= '0';
                    end if;
                elsif(instruction_type = "0010") then
                    if(prime_line_equal_one = '1') then
                        case (operands_size) is
                            when "000" =>
                                -- multiplication_with_reduction_special_prime_0;
                                -- -- In case of size 1
                                -- reg_a = a0_X; reg_b = b0_X; reg_acc = 0; Enable sign a,b; operation : a*b + acc;
                                next_sm_free_flag <= '0';
                                next_sm_rotation_size <= "11";
                                next_sm_circular_shift_enable <= '1';
                                next_sel_address_a <= '0';
                                next_sel_address_b_prime <= "00";
                                next_sm_specific_mac_address_a <= "000";
                                next_sm_specific_mac_address_b <= "000";
                                next_sm_specific_mac_address_o <= "000";
                                next_sm_specific_mac_next_address_o <= "001";
                                next_mac_enable_signed_a <= '0';
                                next_mac_enable_signed_b <= '0';
                                next_mac_sel_load_reg_a <= "00";
                                next_mac_clear_reg_b <= '0';
                                next_mac_clear_reg_acc <= '1';
                                next_mac_sel_shift_reg_o <= '0';
                                next_mac_enable_update_reg_s <= '0';
                                next_mac_sel_reg_s_reg_o_sign <= '0';
                                next_mac_reg_s_reg_o_positive <= '0';
                                next_sm_sign_a_mode <= '0';
                                next_sm_mac_operation_mode <= "10";
                                next_mac_enable_reg_s_mask <= '0';
                                next_mac_subtraction_reg_a_b <= '0';
                                next_mac_sel_multiply_two_a_b <= '0';
                                next_mac_sel_reg_y_output <= '0';
                                next_sm_mac_write_enable_output <= '0';
                                next_mac_memory_double_mode <= '0';
                                next_mac_memory_only_write_mode <= '0';
                                next_base_address_generator_o_increment_previous_address <= '0';
                            when "001"| "010"| "011" =>
                                -- multiplication_with_reduction_special_prime_3;
                                -- -- In case of sizes 2, 3, 4
                                -- reg_a = a0_X; reg_b = b0_X; reg_acc = 0; o0_X = reg_o; operation : a*b + acc;
                                next_sm_free_flag <= '0';
                                next_sm_rotation_size <= "11";
                                next_sm_circular_shift_enable <= '1';
                                next_sel_address_a <= '0';
                                next_sel_address_b_prime <= "00";
                                next_sm_specific_mac_address_a <= "000";
                                next_sm_specific_mac_address_b <= "000";
                                next_sm_specific_mac_address_o <= "000";
                                next_sm_specific_mac_next_address_o <= "001";
                                next_mac_enable_signed_a <= '0';
                                next_mac_enable_signed_b <= '0';
                                next_mac_sel_load_reg_a <= "00";
                                next_mac_clear_reg_b <= '0';
                                next_mac_clear_reg_acc <= '1';
                                next_mac_sel_shift_reg_o <= '0';
                                next_mac_enable_update_reg_s <= '0';
                                next_mac_sel_reg_s_reg_o_sign <= '0';
                                next_mac_reg_s_reg_o_positive <= '0';
                                next_sm_sign_a_mode <= '0';
                                next_sm_mac_operation_mode <= "10";
                                next_mac_enable_reg_s_mask <= '0';
                                next_mac_subtraction_reg_a_b <= '0';
                                next_mac_sel_multiply_two_a_b <= '0';
                                next_mac_sel_reg_y_output <= '0';
                                next_sm_mac_write_enable_output <= '1';
                                next_mac_memory_double_mode <= '0';
                                next_mac_memory_only_write_mode <= '0';
                                next_base_address_generator_o_increment_previous_address <= '0';
                            when "100"| "101" =>
                                -- multiplication_with_reduction_special_prime_47;
                                -- -- In case of sizes 5, 6
                                -- reg_a = a0_X; reg_b = b0_X; reg_acc = 0; o0_X = reg_o; operation : a*b + acc;
                                next_sm_free_flag <= '0';
                                next_sm_rotation_size <= "11";
                                next_sm_circular_shift_enable <= '1';
                                next_sel_address_a <= '0';
                                next_sel_address_b_prime <= "00";
                                next_sm_specific_mac_address_a <= "000";
                                next_sm_specific_mac_address_b <= "000";
                                next_sm_specific_mac_address_o <= "000";
                                next_sm_specific_mac_next_address_o <= "001";
                                next_mac_enable_signed_a <= '0';
                                next_mac_enable_signed_b <= '0';
                                next_mac_sel_load_reg_a <= "00";
                                next_mac_clear_reg_b <= '0';
                                next_mac_clear_reg_acc <= '1';
                                next_mac_sel_shift_reg_o <= '0';
                                next_mac_enable_update_reg_s <= '0';
                                next_mac_sel_reg_s_reg_o_sign <= '0';
                                next_mac_reg_s_reg_o_positive <= '0';
                                next_sm_sign_a_mode <= '0';
                                next_sm_mac_operation_mode <= "10";
                                next_mac_enable_reg_s_mask <= '0';
                                next_mac_subtraction_reg_a_b <= '0';
                                next_mac_sel_multiply_two_a_b <= '0';
                                next_mac_sel_reg_y_output <= '0';
                                next_sm_mac_write_enable_output <= '1';
                                next_mac_memory_double_mode <= '0';
                                next_mac_memory_only_write_mode <= '0';
                                next_base_address_generator_o_increment_previous_address <= '0';
                            when others => 
                                -- multiplication_with_reduction_special_prime_130;
                                -- -- In case of sizes 7, 8
                                -- reg_a = a0_X; reg_b = b0_X; reg_acc = 0; o0_X = reg_o; operation : a*b + acc;
                                next_sm_free_flag <= '0';
                                next_sm_rotation_size <= "11";
                                next_sm_circular_shift_enable <= '1';
                                next_sel_address_a <= '0';
                                next_sel_address_b_prime <= "00";
                                next_sm_specific_mac_address_a <= "000";
                                next_sm_specific_mac_address_b <= "000";
                                next_sm_specific_mac_address_o <= "000";
                                next_sm_specific_mac_next_address_o <= "001";
                                next_mac_enable_signed_a <= '0';
                                next_mac_enable_signed_b <= '0';
                                next_mac_sel_load_reg_a <= "00";
                                next_mac_clear_reg_b <= '0';
                                next_mac_clear_reg_acc <= '1';
                                next_mac_sel_shift_reg_o <= '0';
                                next_mac_enable_update_reg_s <= '0';
                                next_mac_sel_reg_s_reg_o_sign <= '0';
                                next_mac_reg_s_reg_o_positive <= '0';
                                next_sm_sign_a_mode <= '0';
                                next_sm_mac_operation_mode <= "10";
                                next_mac_enable_reg_s_mask <= '0';
                                next_mac_subtraction_reg_a_b <= '0';
                                next_mac_sel_multiply_two_a_b <= '0';
                                next_mac_sel_reg_y_output <= '0';
                                next_sm_mac_write_enable_output <= '1';
                                next_mac_memory_double_mode <= '0';
                                next_mac_memory_only_write_mode <= '0';
                                next_base_address_generator_o_increment_previous_address <= '0';
                        end case;
                    else
                        if(operands_size = "000") then
                            -- multiplication_with_reduction_0;
                            -- -- In case of size 1
                            -- reg_a = a0_X; reg_b = b0_X; reg_acc = 0; Enable sign a,b; operation : a*b + acc;
                            next_sm_free_flag <= '0';
                            next_sm_rotation_size <= "11";
                            next_sm_circular_shift_enable <= '1';
                            next_sel_address_a <= '0';
                            next_sel_address_b_prime <= "00";
                            next_sm_specific_mac_address_a <= "000";
                            next_sm_specific_mac_address_b <= "000";
                            next_sm_specific_mac_address_o <= "000";
                            next_sm_specific_mac_next_address_o <= "001";
                            next_mac_enable_signed_a <= '1';
                            next_mac_enable_signed_b <= '1';
                            next_mac_sel_load_reg_a <= "00";
                            next_mac_clear_reg_b <= '0';
                            next_mac_clear_reg_acc <= '1';
                            next_mac_sel_shift_reg_o <= '0';
                            next_mac_enable_update_reg_s <= '0';
                            next_mac_sel_reg_s_reg_o_sign <= '0';
                            next_mac_reg_s_reg_o_positive <= '0';
                            next_sm_sign_a_mode <= '0';
                            next_sm_mac_operation_mode <= "10";
                            next_mac_enable_reg_s_mask <= '0';
                            next_mac_subtraction_reg_a_b <= '0';
                            next_mac_sel_multiply_two_a_b <= '0';
                            next_mac_sel_reg_y_output <= '0';
                            next_sm_mac_write_enable_output <= '0';
                            next_mac_memory_double_mode <= '0';
                            next_mac_memory_only_write_mode <= '0';
                            next_base_address_generator_o_increment_previous_address <= '0';
                        else
                            -- multiplication_with_reduction_5;
                            -- -- In case of sizes 2, 3, 4, 5, 6, 7, 8
                            -- reg_a = a0_X; reg_b = b0_X; reg_acc = 0; operation : a*b + acc;
                            next_sm_free_flag <= '0';
                            next_sm_rotation_size <= "11";
                            next_sm_circular_shift_enable <= '1';
                            next_sel_address_a <= '0';
                            next_sel_address_b_prime <= "00";
                            next_sm_specific_mac_address_a <= "000";
                            next_sm_specific_mac_address_b <= "000";
                            next_sm_specific_mac_address_o <= "000";
                            next_sm_specific_mac_next_address_o <= "001";
                            next_mac_enable_signed_a <= '0';
                            next_mac_enable_signed_b <= '0';
                            next_mac_sel_load_reg_a <= "00";
                            next_mac_clear_reg_b <= '0';
                            next_mac_clear_reg_acc <= '1';
                            next_mac_sel_shift_reg_o <= '0';
                            next_mac_enable_update_reg_s <= '0';
                            next_mac_sel_reg_s_reg_o_sign <= '0';
                            next_mac_reg_s_reg_o_positive <= '0';
                            next_sm_sign_a_mode <= '0';
                            next_sm_mac_operation_mode <= "10";
                            next_mac_enable_reg_s_mask <= '0';
                            next_mac_subtraction_reg_a_b <= '0';
                            next_mac_sel_multiply_two_a_b <= '0';
                            next_mac_sel_reg_y_output <= '0';
                            next_sm_mac_write_enable_output <= '0';
                            next_mac_memory_double_mode <= '0';
                            next_mac_memory_only_write_mode <= '0';
                            next_base_address_generator_o_increment_previous_address <= '0';
                        end if;
                    end if;
                elsif(instruction_type = "0011") then
                    if(prime_line_equal_one = '1') then
                        case (operands_size) is
                            when "000" =>
                                -- square_with_reduction_special_prime_0;
                                -- -- In case of size 1
                                -- reg_a = a0_X; reg_b = a0_X; reg_acc = 0; Enable sign a,b; operation : a*b + acc;
                                next_sm_free_flag <= '0';
                                next_sm_rotation_size <= "11";
                                next_sm_circular_shift_enable <= '1';
                                next_sel_address_a <= '0';
                                next_sel_address_b_prime <= "00";
                                next_sm_specific_mac_address_a <= "000";
                                next_sm_specific_mac_address_b <= "000";
                                next_sm_specific_mac_address_o <= "000";
                                next_sm_specific_mac_next_address_o <= "001";
                                next_mac_enable_signed_a <= '1';
                                next_mac_enable_signed_b <= '1';
                                next_mac_sel_load_reg_a <= "00";
                                next_mac_clear_reg_b <= '0';
                                next_mac_clear_reg_acc <= '1';
                                next_mac_sel_shift_reg_o <= '0';
                                next_mac_enable_update_reg_s <= '0';
                                next_mac_sel_reg_s_reg_o_sign <= '0';
                                next_mac_reg_s_reg_o_positive <= '0';
                                next_sm_sign_a_mode <= '0';
                                next_sm_mac_operation_mode <= "10";
                                next_mac_enable_reg_s_mask <= '0';
                                next_mac_subtraction_reg_a_b <= '0';
                                next_mac_sel_multiply_two_a_b <= '0';
                                next_mac_sel_reg_y_output <= '0';
                                next_sm_mac_write_enable_output <= '0';
                                next_mac_memory_double_mode <= '0';
                                next_mac_memory_only_write_mode <= '0';
                                next_base_address_generator_o_increment_previous_address <= '0';
                            when "001"| "010"| "011" =>
                                -- square_with_reduction_special_prime_3;
                                -- -- In case of size 2, 3, 4
                                -- reg_a = a0_X; reg_b = a0_X; reg_acc = 0; o0_X = reg_o; operation : a*b + acc;
                                next_sm_free_flag <= '0';
                                next_sm_rotation_size <= "11";
                                next_sm_circular_shift_enable <= '1';
                                next_sel_address_a <= '0';
                                next_sel_address_b_prime <= "00";
                                next_sm_specific_mac_address_a <= "000";
                                next_sm_specific_mac_address_b <= "000";
                                next_sm_specific_mac_address_o <= "000";
                                next_sm_specific_mac_next_address_o <= "001";
                                next_mac_enable_signed_a <= '0';
                                next_mac_enable_signed_b <= '0';
                                next_mac_sel_load_reg_a <= "00";
                                next_mac_clear_reg_b <= '0';
                                next_mac_clear_reg_acc <= '1';
                                next_mac_sel_shift_reg_o <= '0';
                                next_mac_enable_update_reg_s <= '0';
                                next_mac_sel_reg_s_reg_o_sign <= '0';
                                next_mac_reg_s_reg_o_positive <= '0';
                                next_sm_sign_a_mode <= '0';
                                next_sm_mac_operation_mode <= "10";
                                next_mac_enable_reg_s_mask <= '0';
                                next_mac_subtraction_reg_a_b <= '0';
                                next_mac_sel_multiply_two_a_b <= '0';
                                next_mac_sel_reg_y_output <= '0';
                                next_sm_mac_write_enable_output <= '1';
                                next_mac_memory_double_mode <= '0';
                                next_mac_memory_only_write_mode <= '0';
                                next_base_address_generator_o_increment_previous_address <= '0';
                            when "100"| "101" =>
                                -- square_with_reduction_special_prime_37;
                                -- -- In case of size 5, 6
                                -- reg_a = a0_X; reg_b = a0_X; reg_acc = 0; o0_X = reg_o; operation : a*b + acc;
                                next_sm_free_flag <= '0';
                                next_sm_rotation_size <= "11";
                                next_sm_circular_shift_enable <= '1';
                                next_sel_address_a <= '0';
                                next_sel_address_b_prime <= "00";
                                next_sm_specific_mac_address_a <= "000";
                                next_sm_specific_mac_address_b <= "000";
                                next_sm_specific_mac_address_o <= "000";
                                next_sm_specific_mac_next_address_o <= "001";
                                next_mac_enable_signed_a <= '0';
                                next_mac_enable_signed_b <= '0';
                                next_mac_sel_load_reg_a <= "00";
                                next_mac_clear_reg_b <= '0';
                                next_mac_clear_reg_acc <= '1';
                                next_mac_sel_shift_reg_o <= '0';
                                next_mac_enable_update_reg_s <= '0';
                                next_mac_sel_reg_s_reg_o_sign <= '0';
                                next_mac_reg_s_reg_o_positive <= '0';
                                next_sm_sign_a_mode <= '0';
                                next_sm_mac_operation_mode <= "10";
                                next_mac_enable_reg_s_mask <= '0';
                                next_mac_subtraction_reg_a_b <= '0';
                                next_mac_sel_multiply_two_a_b <= '0';
                                next_mac_sel_reg_y_output <= '0';
                                next_sm_mac_write_enable_output <= '1';
                                next_mac_memory_double_mode <= '0';
                                next_mac_memory_only_write_mode <= '0';
                                next_base_address_generator_o_increment_previous_address <= '0';
                            when others => 
                                -- square_with_reduction_special_prime_100;
                                -- -- In case of size 7, 8
                                -- reg_a = a0_X; reg_b = a0_X; reg_acc = 0; o0_X = reg_o; operation : a*b + acc;
                                next_sm_free_flag <= '0';
                                next_sm_rotation_size <= "11";
                                next_sm_circular_shift_enable <= '1';
                                next_sel_address_a <= '0';
                                next_sel_address_b_prime <= "00";
                                next_sm_specific_mac_address_a <= "000";
                                next_sm_specific_mac_address_b <= "000";
                                next_sm_specific_mac_address_o <= "000";
                                next_sm_specific_mac_next_address_o <= "001";
                                next_mac_enable_signed_a <= '0';
                                next_mac_enable_signed_b <= '0';
                                next_mac_sel_load_reg_a <= "00";
                                next_mac_clear_reg_b <= '0';
                                next_mac_clear_reg_acc <= '1';
                                next_mac_sel_shift_reg_o <= '0';
                                next_mac_enable_update_reg_s <= '0';
                                next_mac_sel_reg_s_reg_o_sign <= '0';
                                next_mac_reg_s_reg_o_positive <= '0';
                                next_sm_sign_a_mode <= '0';
                                next_sm_mac_operation_mode <= "10";
                                next_mac_enable_reg_s_mask <= '0';
                                next_mac_subtraction_reg_a_b <= '0';
                                next_mac_sel_multiply_two_a_b <= '0';
                                next_mac_sel_reg_y_output <= '0';
                                next_sm_mac_write_enable_output <= '1';
                                next_mac_memory_double_mode <= '0';
                                next_mac_memory_only_write_mode <= '0';
                                next_base_address_generator_o_increment_previous_address <= '0';
                        end case;
                    else
                        if(operands_size = "000") then
                            -- square_with_reduction_0;
                            -- -- In case of size 1
                            -- reg_a = a0_X; reg_b = a0_X; reg_acc = 0; Enable sign a,b; operation : a*b + acc;
                            next_sm_free_flag <= '0';
                            next_sm_rotation_size <= "11";
                            next_sm_circular_shift_enable <= '1';
                            next_sel_address_a <= '0';
                            next_sel_address_b_prime <= "00";
                            next_sm_specific_mac_address_a <= "000";
                            next_sm_specific_mac_address_b <= "000";
                            next_sm_specific_mac_address_o <= "000";
                            next_sm_specific_mac_next_address_o <= "001";
                            next_mac_enable_signed_a <= '1';
                            next_mac_enable_signed_b <= '1';
                            next_mac_sel_load_reg_a <= "00";
                            next_mac_clear_reg_b <= '0';
                            next_mac_clear_reg_acc <= '1';
                            next_mac_sel_shift_reg_o <= '0';
                            next_mac_enable_update_reg_s <= '0';
                            next_mac_sel_reg_s_reg_o_sign <= '0';
                            next_mac_reg_s_reg_o_positive <= '0';
                            next_sm_sign_a_mode <= '0';
                            next_sm_mac_operation_mode <= "10";
                            next_mac_enable_reg_s_mask <= '0';
                            next_mac_subtraction_reg_a_b <= '0';
                            next_mac_sel_multiply_two_a_b <= '0';
                            next_mac_sel_reg_y_output <= '0';
                            next_sm_mac_write_enable_output <= '0';
                            next_mac_memory_double_mode <= '0';
                            next_mac_memory_only_write_mode <= '0';
                            next_base_address_generator_o_increment_previous_address <= '0';
                        else
                            -- square_with_reduction_5;
                            -- -- In case of 2, 3, 4, 5, 6, 7, 8
                            -- reg_a = a0_X; reg_b = a0_X; reg_acc = 0; operation : a*b + acc;
                            next_sm_free_flag <= '0';
                            next_sm_rotation_size <= "11";
                            next_sm_circular_shift_enable <= '1';
                            next_sel_address_a <= '0';
                            next_sel_address_b_prime <= "00";
                            next_sm_specific_mac_address_a <= "000";
                            next_sm_specific_mac_address_b <= "000";
                            next_sm_specific_mac_address_o <= "000";
                            next_sm_specific_mac_next_address_o <= "001";
                            next_mac_enable_signed_a <= '0';
                            next_mac_enable_signed_b <= '0';
                            next_mac_sel_load_reg_a <= "00";
                            next_mac_clear_reg_b <= '0';
                            next_mac_clear_reg_acc <= '1';
                            next_mac_sel_shift_reg_o <= '0';
                            next_mac_enable_update_reg_s <= '0';
                            next_mac_sel_reg_s_reg_o_sign <= '0';
                            next_mac_reg_s_reg_o_positive <= '0';
                            next_sm_sign_a_mode <= '0';
                            next_sm_mac_operation_mode <= "10";
                            next_mac_enable_reg_s_mask <= '0';
                            next_mac_subtraction_reg_a_b <= '0';
                            next_mac_sel_multiply_two_a_b <= '0';
                            next_mac_sel_reg_y_output <= '0';
                            next_sm_mac_write_enable_output <= '0';
                            next_mac_memory_double_mode <= '0';
                            next_mac_memory_only_write_mode <= '0';
                            next_base_address_generator_o_increment_previous_address <= '0';
                        end if;
                    end if;
                elsif(instruction_type = "0100") then
                    if(operands_size = "000") then
                        -- addition_subtraction_direct_0;
                        -- -- In case of size 1
                        -- reg_a = a0_X; reg_b = b0_X; reg_acc = 0; o0_0 = reg_o; Enable sign a,b; operation : b +/- a + acc;
                        next_sm_free_flag <= '0';
                        next_sm_rotation_size <= "10";
                        next_sm_circular_shift_enable <= '1';
                        next_sel_address_a <= '0';
                        next_sel_address_b_prime <= "00";
                        next_sm_specific_mac_address_a <= "000";
                        next_sm_specific_mac_address_b <= "000";
                        next_sm_specific_mac_address_o <= "000";
                        next_sm_specific_mac_next_address_o <= "001";
                        next_mac_enable_signed_a <= '1';
                        next_mac_enable_signed_b <= '1';
                        next_mac_sel_load_reg_a <= "00";
                        next_mac_clear_reg_b <= '0';
                        next_mac_clear_reg_acc <= '1';
                        next_mac_sel_shift_reg_o <= '0';
                        next_mac_enable_update_reg_s <= '0';
                        next_mac_sel_reg_s_reg_o_sign <= '0';
                        next_mac_reg_s_reg_o_positive <= '0';
                        next_sm_sign_a_mode <= '1';
                        next_sm_mac_operation_mode(1) <= '0';
                        next_sm_mac_operation_mode(0) <= '0';
                        next_mac_enable_reg_s_mask <= '0';
                        next_mac_subtraction_reg_a_b <= '0';
                        next_mac_sel_multiply_two_a_b <= '0';
                        next_mac_sel_reg_y_output <= '0';
                        next_sm_mac_write_enable_output <= '1';
                        next_mac_memory_double_mode <= '0';
                        next_mac_memory_only_write_mode <= '0';
                        next_base_address_generator_o_increment_previous_address <= '0';
                    else
                        -- addition_subtraction_direct_2;
                        -- -- In case of size 2, 3, 4, 5, 6, 7, 8
                        -- reg_a = a0_X; reg_b = b0_X; reg_acc = 0; o0_X = reg_o; operation : b +/- a + acc;
                        next_sm_free_flag <= '0';
                        next_sm_rotation_size <= "10";
                        next_sm_circular_shift_enable <= '1';
                        next_sel_address_a <= '0';
                        next_sel_address_b_prime <= "00";
                        next_sm_specific_mac_address_a <= "000";
                        next_sm_specific_mac_address_b <= "000";
                        next_sm_specific_mac_address_o <= "000";
                        next_sm_specific_mac_next_address_o <= "001";
                        next_mac_enable_signed_a <= '0';
                        next_mac_enable_signed_b <= '0';
                        next_mac_sel_load_reg_a <= "00";
                        next_mac_clear_reg_b <= '0';
                        next_mac_clear_reg_acc <= '1';
                        next_mac_sel_shift_reg_o <= '0';
                        next_mac_enable_update_reg_s <= '0';
                        next_mac_sel_reg_s_reg_o_sign <= '0';
                        next_mac_reg_s_reg_o_positive <= '0';
                        next_sm_sign_a_mode <= '1';
                        next_sm_mac_operation_mode(1) <= '0';
                        next_sm_mac_operation_mode(0) <= '0';
                        next_mac_enable_reg_s_mask <= '0';
                        next_mac_subtraction_reg_a_b <= '0';
                        next_mac_sel_multiply_two_a_b <= '0';
                        next_mac_sel_reg_y_output <= '0';
                        next_sm_mac_write_enable_output <= '1';
                        next_mac_memory_double_mode <= '0';
                        next_mac_memory_only_write_mode <= '0';
                        next_base_address_generator_o_increment_previous_address <= '0';
                    end if;
                elsif(instruction_type = "0101") then
                    if(operands_size = "000") then
                        -- iterative_modular_reduction_0;
                        -- -- In case of size 1
                        -- reg_a = a0_X; reg_b = 0; reg_acc = 0; Enable sign a,b; operation : b + a + acc;
                        next_sm_free_flag <= '0';
                        next_sm_rotation_size <= "10";
                        next_sm_circular_shift_enable <= '1';
                        next_sel_address_a <= '0';
                        next_sel_address_b_prime <= "10";
                        next_sm_specific_mac_address_a <= "000";
                        next_sm_specific_mac_address_b <= "000";
                        next_sm_specific_mac_address_o <= "000";
                        next_sm_specific_mac_next_address_o <= "001";
                        next_mac_enable_signed_a <= '1';
                        next_mac_enable_signed_b <= '1';
                        next_mac_sel_load_reg_a <= "00";
                        next_mac_clear_reg_b <= '1';
                        next_mac_clear_reg_acc <= '1';
                        next_mac_sel_shift_reg_o <= '0';
                        next_mac_enable_update_reg_s <= '0';
                        next_mac_sel_reg_s_reg_o_sign <= '0';
                        next_mac_reg_s_reg_o_positive <= '0';
                        next_sm_sign_a_mode <= '0';
                        next_sm_mac_operation_mode <= "01";
                        next_mac_enable_reg_s_mask <= '0';
                        next_mac_subtraction_reg_a_b <= '0';
                        next_mac_sel_multiply_two_a_b <= '0';
                        next_mac_sel_reg_y_output <= '0';
                        next_sm_mac_write_enable_output <= '0';
                        next_mac_memory_double_mode <= '0';
                        next_mac_memory_only_write_mode <= '0';
                        next_base_address_generator_o_increment_previous_address <= '0';
                    elsif(operands_size = "001") then
                        -- iterative_modular_reduction_5;
                        -- -- In case of size 2
                        -- reg_a = a1_X; reg_b = 0; reg_acc = 0; Enable sign a,b; operation : b + a + acc;
                        next_sm_free_flag <= '0';
                        next_sm_rotation_size <= "10";
                        next_sm_circular_shift_enable <= '1';
                        next_sel_address_a <= '0';
                        next_sel_address_b_prime <= "10";
                        next_sm_specific_mac_address_a <= "001";
                        next_sm_specific_mac_address_b <= "000";
                        next_sm_specific_mac_address_o <= "000";
                        next_sm_specific_mac_next_address_o <= "001";
                        next_mac_enable_signed_a <= '1';
                        next_mac_enable_signed_b <= '1';
                        next_mac_sel_load_reg_a <= "00";
                        next_mac_clear_reg_b <= '1';
                        next_mac_clear_reg_acc <= '1';
                        next_mac_sel_shift_reg_o <= '0';
                        next_mac_enable_update_reg_s <= '0';
                        next_mac_sel_reg_s_reg_o_sign <= '0';
                        next_mac_reg_s_reg_o_positive <= '0';
                        next_sm_sign_a_mode <= '0';
                        next_sm_mac_operation_mode <= "01";
                        next_mac_enable_reg_s_mask <= '0';
                        next_mac_subtraction_reg_a_b <= '0';
                        next_mac_sel_multiply_two_a_b <= '0';
                        next_mac_sel_reg_y_output <= '0';
                        next_sm_mac_write_enable_output <= '0';
                        next_mac_memory_double_mode <= '0';
                        next_mac_memory_only_write_mode <= '0';
                        next_base_address_generator_o_increment_previous_address <= '0';
                    elsif(operands_size = "010") then
                        -- iterative_modular_reduction_13;
                        -- -- In case of size 3
                        -- reg_a = a2_X; reg_b = 0; reg_acc = 0; Enable sign a,b; operation : b + a + acc;
                        next_sm_free_flag <= '0';
                        next_sm_rotation_size <= "10";
                        next_sm_circular_shift_enable <= '1';
                        next_sel_address_a <= '0';
                        next_sel_address_b_prime <= "10";
                        next_sm_specific_mac_address_a <= "010";
                        next_sm_specific_mac_address_b <= "010";
                        next_sm_specific_mac_address_o <= "010";
                        next_sm_specific_mac_next_address_o <= "011";
                        next_mac_enable_signed_a <= '1';
                        next_mac_enable_signed_b <= '1';
                        next_mac_sel_load_reg_a <= "00";
                        next_mac_clear_reg_b <= '1';
                        next_mac_clear_reg_acc <= '1';
                        next_mac_sel_shift_reg_o <= '0';
                        next_mac_enable_update_reg_s <= '0';
                        next_mac_sel_reg_s_reg_o_sign <= '0';
                        next_mac_reg_s_reg_o_positive <= '0';
                        next_sm_sign_a_mode <= '0';
                        next_sm_mac_operation_mode <= "01";
                        next_mac_enable_reg_s_mask <= '0';
                        next_mac_subtraction_reg_a_b <= '0';
                        next_mac_sel_multiply_two_a_b <= '0';
                        next_mac_sel_reg_y_output <= '0';
                        next_sm_mac_write_enable_output <= '0';
                        next_mac_memory_double_mode <= '0';
                        next_mac_memory_only_write_mode <= '0';
                        next_base_address_generator_o_increment_previous_address <= '0';
                    elsif(operands_size = "011") then
                        -- iterative_modular_reduction_24;
                        -- -- In case of size 4
                        -- reg_a = a3_X; reg_b = 0; reg_acc = 0; Enable sign a,b; operation : b + a + acc;
                        next_sm_free_flag <= '0';
                        next_sm_rotation_size <= "10";
                        next_sm_circular_shift_enable <= '1';
                        next_sel_address_a <= '0';
                        next_sel_address_b_prime <= "10";
                        next_sm_specific_mac_address_a <= "011";
                        next_sm_specific_mac_address_b <= "011";
                        next_sm_specific_mac_address_o <= "011";
                        next_sm_specific_mac_next_address_o <= "000";
                        next_mac_enable_signed_a <= '1';
                        next_mac_enable_signed_b <= '1';
                        next_mac_sel_load_reg_a <= "00";
                        next_mac_clear_reg_b <= '1';
                        next_mac_clear_reg_acc <= '1';
                        next_mac_sel_shift_reg_o <= '0';
                        next_mac_enable_update_reg_s <= '0';
                        next_mac_sel_reg_s_reg_o_sign <= '0';
                        next_mac_reg_s_reg_o_positive <= '0';
                        next_sm_sign_a_mode <= '0';
                        next_sm_mac_operation_mode <= "01";
                        next_mac_enable_reg_s_mask <= '0';
                        next_mac_subtraction_reg_a_b <= '0';
                        next_mac_sel_multiply_two_a_b <= '0';
                        next_mac_sel_reg_y_output <= '0';
                        next_sm_mac_write_enable_output <= '0';
                        next_mac_memory_double_mode <= '0';
                        next_mac_memory_only_write_mode <= '0';
                        next_base_address_generator_o_increment_previous_address <= '0';
                    elsif(operands_size = "100") then
                        -- iterative_modular_reduction_38;
                        -- -- In case of size 5
                        -- reg_a = a4_X; reg_b = 0; reg_acc = 0; Enable sign a,b; operation : b + a + acc;
                        next_sm_free_flag <= '0';
                        next_sm_rotation_size <= "10";
                        next_sm_circular_shift_enable <= '1';
                        next_sel_address_a <= '0';
                        next_sel_address_b_prime <= "10";
                        next_sm_specific_mac_address_a <= "100";
                        next_sm_specific_mac_address_b <= "100";
                        next_sm_specific_mac_address_o <= "100";
                        next_sm_specific_mac_next_address_o <= "101";
                        next_mac_enable_signed_a <= '1';
                        next_mac_enable_signed_b <= '1';
                        next_mac_sel_load_reg_a <= "00";
                        next_mac_clear_reg_b <= '1';
                        next_mac_clear_reg_acc <= '1';
                        next_mac_sel_shift_reg_o <= '0';
                        next_mac_enable_update_reg_s <= '0';
                        next_mac_sel_reg_s_reg_o_sign <= '0';
                        next_mac_reg_s_reg_o_positive <= '0';
                        next_sm_sign_a_mode <= '0';
                        next_sm_mac_operation_mode <= "01";
                        next_mac_enable_reg_s_mask <= '0';
                        next_mac_subtraction_reg_a_b <= '0';
                        next_mac_sel_multiply_two_a_b <= '0';
                        next_mac_sel_reg_y_output <= '0';
                        next_sm_mac_write_enable_output <= '0';
                        next_mac_memory_double_mode <= '0';
                        next_mac_memory_only_write_mode <= '0';
                        next_base_address_generator_o_increment_previous_address <= '0';
                    elsif(operands_size = "101") then
                        -- iterative_modular_reduction_55;
                        -- -- In case of size 6
                        -- reg_a = a5_X; reg_b = 0; reg_acc = 0; Enable sign a,b; operation : b + a + acc;
                        next_sm_free_flag <= '0';
                        next_sm_rotation_size <= "10";
                        next_sm_circular_shift_enable <= '1';
                        next_sel_address_a <= '0';
                        next_sel_address_b_prime <= "10";
                        next_sm_specific_mac_address_a <= "101";
                        next_sm_specific_mac_address_b <= "101";
                        next_sm_specific_mac_address_o <= "101";
                        next_sm_specific_mac_next_address_o <= "110";
                        next_mac_enable_signed_a <= '1';
                        next_mac_enable_signed_b <= '1';
                        next_mac_sel_load_reg_a <= "00";
                        next_mac_clear_reg_b <= '1';
                        next_mac_clear_reg_acc <= '1';
                        next_mac_sel_shift_reg_o <= '0';
                        next_mac_enable_update_reg_s <= '0';
                        next_mac_sel_reg_s_reg_o_sign <= '0';
                        next_mac_reg_s_reg_o_positive <= '0';
                        next_sm_sign_a_mode <= '0';
                        next_sm_mac_operation_mode <= "01";
                        next_mac_enable_reg_s_mask <= '0';
                        next_mac_subtraction_reg_a_b <= '0';
                        next_mac_sel_multiply_two_a_b <= '0';
                        next_mac_sel_reg_y_output <= '0';
                        next_sm_mac_write_enable_output <= '0';
                        next_mac_memory_double_mode <= '0';
                        next_mac_memory_only_write_mode <= '0';
                        next_base_address_generator_o_increment_previous_address <= '0';
                    elsif(operands_size = "110") then
                        -- iterative_modular_reduction_75;
                        -- -- In case of size 7
                        -- reg_a = a6_X; reg_b = 0; reg_acc = 0; Enable sign a,b; operation : b + a + acc;
                        next_sm_free_flag <= '0';
                        next_sm_rotation_size <= "10";
                        next_sm_circular_shift_enable <= '1';
                        next_sel_address_a <= '0';
                        next_sel_address_b_prime <= "10";
                        next_sm_specific_mac_address_a <= "110";
                        next_sm_specific_mac_address_b <= "110";
                        next_sm_specific_mac_address_o <= "110";
                        next_sm_specific_mac_next_address_o <= "111";
                        next_mac_enable_signed_a <= '1';
                        next_mac_enable_signed_b <= '1';
                        next_mac_sel_load_reg_a <= "00";
                        next_mac_clear_reg_b <= '1';
                        next_mac_clear_reg_acc <= '1';
                        next_mac_sel_shift_reg_o <= '0';
                        next_mac_enable_update_reg_s <= '0';
                        next_mac_sel_reg_s_reg_o_sign <= '0';
                        next_mac_reg_s_reg_o_positive <= '0';
                        next_sm_sign_a_mode <= '0';
                        next_sm_mac_operation_mode <= "01";
                        next_mac_enable_reg_s_mask <= '0';
                        next_mac_subtraction_reg_a_b <= '0';
                        next_mac_sel_multiply_two_a_b <= '0';
                        next_mac_sel_reg_y_output <= '0';
                        next_sm_mac_write_enable_output <= '0';
                        next_mac_memory_double_mode <= '0';
                        next_mac_memory_only_write_mode <= '0';
                        next_base_address_generator_o_increment_previous_address <= '0';
                    else
                        -- iterative_modular_reduction_98;
                        -- -- In case of size 8
                        -- reg_a = a7_X; reg_b = 0; reg_acc = 0; Enable sign a,b; operation : b + a + acc;
                        next_sm_free_flag <= '0';
                        next_sm_rotation_size <= "10";
                        next_sm_circular_shift_enable <= '1';
                        next_sel_address_a <= '0';
                        next_sel_address_b_prime <= "10";
                        next_sm_specific_mac_address_a <= "111";
                        next_sm_specific_mac_address_b <= "111";
                        next_sm_specific_mac_address_o <= "111";
                        next_sm_specific_mac_next_address_o <= "000";
                        next_mac_enable_signed_a <= '1';
                        next_mac_enable_signed_b <= '1';
                        next_mac_sel_load_reg_a <= "00";
                        next_mac_clear_reg_b <= '1';
                        next_mac_clear_reg_acc <= '1';
                        next_mac_sel_shift_reg_o <= '0';
                        next_mac_enable_update_reg_s <= '0';
                        next_mac_sel_reg_s_reg_o_sign <= '0';
                        next_mac_reg_s_reg_o_positive <= '0';
                        next_sm_sign_a_mode <= '0';
                        next_sm_mac_operation_mode <= "01";
                        next_mac_enable_reg_s_mask <= '0';
                        next_mac_subtraction_reg_a_b <= '0';
                        next_mac_sel_multiply_two_a_b <= '0';
                        next_mac_sel_reg_y_output <= '0';
                        next_sm_mac_write_enable_output <= '0';
                        next_mac_memory_double_mode <= '0';
                        next_mac_memory_only_write_mode <= '0';
                        next_base_address_generator_o_increment_previous_address <= '0';
                    end if;
                end if;
            end if;
        when multiplication_direct_0 =>
            -- -- In case of size 1
            -- reg_a = a0_X; reg_b = b0_X; reg_acc = 0; o0_X = reg_o; o1_X = reg_o >> 272; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_2 =>
            -- -- Other cases
            -- reg_a = a0_X; reg_b = b0_X; reg_acc = 0; o0_X = reg_o; operation : a*b + acc; o0_X = reg_o;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_3 =>
            -- -- In case of size 2
            -- reg_a = a1_X; reg_b = b0_X; reg_acc = reg_o >> 272; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_4 =>
            -- reg_a = a0_X; reg_b = b1_X; reg_acc = reg_o; o1_X = reg_o; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_5 =>
            -- reg_a = a1_X; reg_b = b1_X; reg_acc = reg_o >> 272; o2_X = reg_o; o3_X = reg_o >> 272; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_7 =>
            -- -- Other cases
            -- reg_a = a1_X; reg_b = b0_X; reg_acc = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_8 =>
            -- reg_a = a0_X; reg_b = b1_X; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_9 =>
            -- reg_a = a1_X; reg_b = b1_X; reg_acc = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_10 =>
            -- -- In case of size 3
            -- reg_a = a0_X; reg_b = b2_X; reg_acc = reg_o; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_11 =>
            -- reg_a = a2_X; reg_b = b0_X; reg_acc = reg_o; Enable sign a; o2_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_12 =>
            -- reg_a = a2_X; reg_b = b1_X; reg_acc = reg_o >> 272; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_13 =>
            -- reg_a = a1_X; reg_b = b2_X; reg_acc = reg_o; o3_X = reg_o; Enable sign b; operation : a*b + acc; 
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_14 =>
            -- reg_a = a2_X; reg_b = b2_X; reg_acc = reg_o >> 272; o4_X = reg_o; o5_X = reg_o >> 272; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_16 =>
            -- -- Other cases
            -- reg_a = a0_0; reg_b = b2_0; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_17 =>
            -- reg_a = a2_X; reg_b = b0_X; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_18 =>
            -- reg_a = a2_X; reg_b = b1_X; reg_acc = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_19 =>
            -- reg_a = a1_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc; 
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_20 =>
            -- -- In case of size 4
            -- reg_a = a3_X; reg_b = b0_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_21 =>
            -- reg_a = a0_X; reg_b = b3_X; reg_acc = reg_o; o3_X = reg_o; Enable sign b; operation : a*b + acc; 
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_22 =>
            -- reg_a = a2_X; reg_b = b2_X; reg_acc = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_23 =>
            -- reg_a = a3_X; reg_b = b1_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_24 =>
            -- reg_a = a1_X; reg_b = b3_X; reg_acc = reg_o; o4_X = reg_o; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_25 =>
            -- reg_a = a3_X; reg_b = b2_X; reg_acc = reg_o >> 272; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_26 =>
            -- reg_a = a2_X; reg_b = b3_X; reg_acc = reg_o; o5_X = reg_o; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_27 =>
            -- reg_a = a3_X; reg_b = b3_X; reg_acc = reg_o >> 272; o6_X = reg_o; o7_X = reg_o >> 272; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_29 =>
            -- -- Other cases
            -- reg_a = a3_X; reg_b = b0_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_30 =>
            -- reg_a = a0_X; reg_b = b3_X; reg_acc = reg_o; o3_0 = reg_o; operation : a*b + acc; 
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_31 =>
            -- reg_a = a2_X; reg_b = b2_X; reg_acc = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_32 =>
            -- reg_a = a3_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_33 =>
            -- reg_a = a1_X; reg_b = b3_X; reg_acc = reg_o; o4_0 = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_34 =>
            -- -- In case of size 5
            -- reg_a = a4_X; reg_b = b0_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_35 =>
            -- reg_a = a0_X; reg_b = b4_X; reg_acc = reg_o; o4_0 = reg_o; Enable sign b; operation : a*b + acc; 
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_36 =>
            -- reg_a = a3_X; reg_b = b2_X; reg_acc = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_37 =>
            -- reg_a = a2_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_38 =>
            -- reg_a = a4_X; reg_b = b1_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_39 =>
            -- reg_a = a1_X; reg_b = b4_X; reg_acc = reg_o; o5_X = reg_o; Enable sign b; operation : a*b + acc; 
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_40 =>
            -- reg_a = a3_X; reg_b = b3_X; reg_acc = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_41 =>
            -- reg_a = a4_X; reg_b = b2_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_42 =>
            -- reg_a = a2_X; reg_b = b4_X; reg_acc = reg_o; o6_X = reg_o; Enable sign b; operation : a*b + acc; 
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_43 =>
            -- reg_a = a4_X; reg_b = b3_X; reg_acc = reg_o >> 272; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "111";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_44 =>
            -- reg_a = a3_X; reg_b = b4_X; reg_acc = reg_o; o7_X = reg_o; Enable sign b; operation : a*b + acc; Increment base address o;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "111";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '1';
        when multiplication_direct_45 =>
            -- reg_a = a4_X; reg_b = b4_X; reg_acc = reg_o >> 272; o8_X = reg_o; o9_X = reg_o >> 272; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_47 =>
            -- -- Other cases
            -- reg_a = a4_X; reg_b = b0_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_48 =>
            -- reg_a = a0_X; reg_b = b4_X; reg_acc = reg_o; o4_X = reg_o; operation : a*b + acc; 
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_49 =>
            -- reg_a = a3_X; reg_b = b2_X; reg_acc = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_50 =>
            -- reg_a = a2_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_51 =>
            -- reg_a = a4_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_52 =>
            -- reg_a = a1_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc; 
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_53 =>
            -- -- In case of size 6
            -- reg_a = a5_X; reg_b = b0_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_54 =>
            -- reg_a = a0_X; reg_b = b5_X; reg_acc = reg_o; o5_0 = reg_o; Enable sign b; operation : a*b + acc; 
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_55 =>
            -- reg_a = a3_X; reg_b = b3_X; reg_acc = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_56 =>
            -- reg_a = a2_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_57 =>
            -- reg_a = a4_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_58 =>
            -- reg_a = a5_X; reg_b = b1_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_59 =>
            -- reg_a = a1_X; reg_b = b5_X; reg_acc = reg_o; o6_0 = reg_o; Enable sign b; operation : a*b + acc; 
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_60 =>
            -- reg_a = a4_X; reg_b = b3_X; reg_acc = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "111";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_61 =>
            -- reg_a = a3_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "111";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_62 =>
            -- reg_a = a5_X; reg_b = b2_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "111";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_63 =>
            -- reg_a = a2_X; reg_b = b5_X; reg_acc = reg_o; o7_0 = reg_o; Enable sign b; operation : a*b + acc; Increment base address o;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "111";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '1';
        when multiplication_direct_64 =>
            -- reg_a = a4_X; reg_b = b4_X; reg_acc = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_65 =>
            -- reg_a = a5_X; reg_b = b3_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_66 =>
            -- reg_a = a3_X; reg_b = b5_X; reg_acc = reg_o; o8_0 = reg_o; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_67 =>
            -- reg_a = a5_X; reg_b = b4_X; reg_acc = reg_o >> 272; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_68 =>
            -- reg_a = a4_X; reg_b = b5_X; reg_acc = reg_o; o9_0 = reg_o; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_69 =>
            -- reg_a = a5_X; reg_b = b5_X; reg_acc = reg_o >> 272; o10_X = reg_o; o11_X = reg_o >> 272; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_71 =>
            -- -- Other cases
            -- reg_a = a5_X; reg_b = b0_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_72 =>
            -- reg_a = a0_X; reg_b = b5_X; reg_acc = reg_o; o5_0 = reg_o; operation : a*b + acc; 
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_73 =>
            -- reg_a = a3_X; reg_b = b3_X; reg_acc = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_74 =>
            -- reg_a = a4_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_75 =>
            -- reg_a = a2_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_76 =>
            -- reg_a = a5_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_77 =>
            -- reg_a = a1_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_78 =>
            -- -- In case of size 7
            -- reg_a = a6_X; reg_b = b0_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_79 =>
            -- reg_a = a0_X; reg_b = b6_X; reg_acc = reg_o; o6_0 = reg_o; Enable sign b; operation : a*b + acc; 
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_80 =>
            -- reg_a = a4_X; reg_b = b3_X; reg_acc = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "111";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_81 =>
            -- reg_a = a3_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "111";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_82 =>
            -- reg_a = a5_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "111";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_83 =>
            -- reg_a = a2_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "111";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_84 =>
            -- reg_a = a6_X; reg_b = b1_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "111";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_85 =>
            -- reg_a = a1_X; reg_b = b6_X; reg_acc = reg_o; o7_0 = reg_o; Enable sign b; operation : a*b + acc; Increment base address o;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "111";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '1';
        when multiplication_direct_86 =>
            -- reg_a = a4_X; reg_b = b4_X; reg_acc = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_87 =>
            -- reg_a = a5_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_88 =>
            -- reg_a = a3_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_89 =>
            -- reg_a = a6_X; reg_b = b2_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_90 =>
            -- reg_a = a2_X; reg_b = b6_X; reg_acc = reg_o; o8_0 = reg_o; Enable sign b; operation : a*b + acc; 
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_91 =>
            -- reg_a = a5_X; reg_b = b4_X; reg_acc = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_92 =>
            -- reg_a = a4_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_93 =>
            -- reg_a = a6_X; reg_b = b3_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_94 =>
            -- reg_a = a3_X; reg_b = b6_X; reg_acc = reg_o; o9_0 = reg_o; Enable sign b; operation : a*b + acc; 
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_95 =>
            -- reg_a = a5_X; reg_b = b5_X; reg_acc = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_96 =>
            -- reg_a = a6_X; reg_b = b4_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_97 =>
            -- reg_a = a4_X; reg_b = b6_X; reg_acc = reg_o; o10_0 = reg_o; Enable sign b; operation : a*b + acc; 
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_98 =>
            -- reg_a = a6_X; reg_b = b5_X; reg_acc = reg_o >> 272; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_99 =>
            -- reg_a = a5_X; reg_b = b6_X; reg_acc = reg_o; o11_0 = reg_o; Enable sign b; operation : a*b + acc; 
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_100 =>
            -- reg_a = a6_X; reg_b = b6_X; reg_acc = reg_o >> 272; o12_X = reg_o; o13_X = reg_o >> 272; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_102 =>
            -- -- In case of size 8
            -- reg_a = a6_X; reg_b = b0_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_103 =>
            -- reg_a = a0_X; reg_b = b6_X; reg_acc = reg_o; o6_0 = reg_o; operation : a*b + acc; 
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_104 =>
            -- reg_a = a4_X; reg_b = b3_X; reg_acc = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "111";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_105 =>
            -- reg_a = a3_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "111";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_106 =>
            -- reg_a = a5_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "111";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_107 =>
            -- reg_a = a2_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "111";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_108 =>
            -- reg_a = a6_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "111";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_109 =>
            -- reg_a = a1_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "111";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_110 =>
            -- reg_a = a7_X; reg_b = b0_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "111";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_111 =>
            -- reg_a = a0_X; reg_b = b7_X; reg_acc = reg_o; o7_0 = reg_o; Enable sign b; operation : a*b + acc; Increment base address o;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "111";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '1';
        when multiplication_direct_112 =>
            -- reg_a = a4_X; reg_b = b4_X; reg_acc = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_113 =>
            -- reg_a = a5_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_114 =>
            -- reg_a = a3_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_115 =>
            -- reg_a = a6_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_116 =>
            -- reg_a = a2_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_117 =>
            -- reg_a = a7_X; reg_b = b1_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_118 =>
            -- reg_a = a1_X; reg_b = b7_X; reg_acc = reg_o; o8_0 = reg_o; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_119 =>
            -- reg_a = a5_X; reg_b = b4_X; reg_acc = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_120 =>
            -- reg_a = a4_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_121 =>
            -- reg_a = a6_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_122 =>
            -- reg_a = a3_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_123 =>
            -- reg_a = a7_X; reg_b = b2_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_124 =>
            -- reg_a = a2_X; reg_b = b7_X; reg_acc = reg_o; o9_0 = reg_o; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_125 =>
            -- reg_a = a5_X; reg_b = b5_X; reg_acc = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_126 =>
            -- reg_a = a6_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_127 =>
            -- reg_a = a4_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_128 =>
            -- reg_a = a7_X; reg_b = b3_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_129 =>
            -- reg_a = a3_X; reg_b = b7_X; reg_acc = reg_o; o10_0 = reg_o; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_130 =>
            -- reg_a = a6_X; reg_b = b5_X; reg_acc = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_131 =>
            -- reg_a = a5_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_132 =>
            -- reg_a = a7_X; reg_b = b4_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_133 =>
            -- reg_a = a4_X; reg_b = b7_X; reg_acc = reg_o; o11_0 = reg_o; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_134 =>
            -- reg_a = a6_X; reg_b = b6_X; reg_acc = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_135 =>
            -- reg_a = a7_X; reg_b = b5_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_136 =>
            -- reg_a = a5_X; reg_b = b7_X; reg_acc = reg_o; o12_0 = reg_o; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_137 =>
            -- reg_a = a7_X; reg_b = b6_X; reg_acc = reg_o >> 272; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_138 =>
            -- reg_a = a6_X; reg_b = b7_X; reg_acc = reg_o; o13_0 = reg_o; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_139 =>
            -- reg_a = a7_X; reg_b = b7_X; reg_acc = reg_o >> 272; o14_X = reg_o; o15_X = reg_o >> 272; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_0 => 
            -- -- In case of size 1
            -- reg_a = a0_X; reg_b = a0_X; reg_acc = 0; o0_X = reg_o; o1_X = reg_o >> 272; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_2 => 
            -- -- In case of sizes 2, 3, 4, 5, 6, 7, 8
            -- reg_a = a0_X; reg_b = a0_X; reg_acc = 0; o0_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_3 => 
            -- -- In case of size 2
            -- reg_a = a1_X; reg_b = a0_X; reg_acc = reg_o >> 272; o1_X = reg_o; Enable sign a; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_4 => 
            -- reg_a = a1_X; reg_b = a1_X; reg_acc = reg_o >> 272; o2_X = reg_o; o3_X = reg_o >> 272; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_6 => 
            -- -- Other cases
            -- reg_a = a1_X; reg_b = a0_X; reg_acc = reg_o >> 272; o1_X = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_7 =>
            -- reg_a = a1_X; reg_b = a1_X; reg_acc = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_8 =>
            -- -- In case of size 3
            -- reg_a = a0_X; reg_b = a2_X; reg_acc = reg_o; o2_X = reg_o; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_9 =>
            -- reg_a = a2_X; reg_b = a1_X; reg_acc = reg_o >> 272; o3_X = reg_o; Enable sign a; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_10 =>
            -- reg_a = a2_X; reg_b = a2_X; reg_acc = reg_o >> 272; o4_X = reg_o; o5_X = reg_o >> 272; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_12 =>
            -- -- Other cases
            -- reg_a = a0_X; reg_b = a2_X; reg_acc = reg_o; o2_X = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_13 =>
            -- reg_a = a2_X; reg_b = a1_X; reg_acc = reg_o >> 272; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_14 =>
            -- -- In case of size 4
            -- reg_a = a3_X; reg_b = a0_X; reg_acc = reg_o; o3_X = reg_o; Enable sign a; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_15 =>
            -- reg_a = a2_X; reg_b = a2_X; reg_acc = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_16 =>
            -- reg_a = a3_X; reg_b = a1_X; reg_acc = reg_o; o4_X = reg_o; Enable sign a; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_17 =>
            -- reg_a = a3_X; reg_b = a2_X; reg_acc = reg_o >> 272; o5_X = reg_o; Enable sign a; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_18 =>
            -- reg_a = a3_X; reg_b = a3_X; reg_acc = reg_o >> 272; o6_X = reg_o; o7_X = reg_o >> 272; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_20 =>
            -- -- Other cases
            -- reg_a = a3_X; reg_b = a0_X; reg_acc = reg_o; o3_X = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_21 =>
            -- reg_a = a2_X; reg_b = a2_X; reg_acc = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_22 =>
            -- reg_a = a3_X; reg_b = a1_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_23 =>
            -- -- In case of size 5
            -- reg_a = a4_X; reg_b = a0_X; reg_acc = reg_o; o4_X = reg_o; Enable sign a; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_24 =>
            -- reg_a = a3_X; reg_b = a2_X; reg_acc = reg_o >> 272; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_25 =>
            -- reg_a = a4_X; reg_b = a1_X; reg_acc = reg_o; o5_X = reg_o; Enable sign a; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_26 =>
            -- reg_a = a3_X; reg_b = a3_X; reg_acc = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_27 =>
            -- reg_a = a4_X; reg_b = a2_X; reg_acc = reg_o; o6_X = reg_o; Enable sign a; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_28 =>
            -- reg_a = a4_X; reg_b = a3_X; reg_acc = reg_o >> 272; o7_X = reg_o; Enable sign a; operation : 2*a*b + acc; Increase base address o;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "111";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '1';
        when square_direct_29 =>
            -- reg_a = a4_X; reg_b = a4_X; reg_acc = reg_o >> 272; o8_X = reg_o; o9_X = reg_o >> 272; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_31 =>
            -- -- Other cases
            -- reg_a = a4_X; reg_b = a0_X; reg_acc = reg_o; o4_X = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_32 =>
            -- reg_a = a3_X; reg_b = a2_X; reg_acc = reg_o >> 272; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_33 =>
            -- reg_a = a4_X; reg_b = a1_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_34 =>
            -- -- In case of size 6
            -- reg_a = a5_X; reg_b = a0_X; reg_acc = reg_o; o5_X = reg_o; Enable sign a; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_35 =>
            -- reg_a = a3_X; reg_b = a3_X; reg_acc = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_36 =>
            -- reg_a = a4_X; reg_b = a2_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_37 =>
            -- reg_a = a5_X; reg_b = a1_X; reg_acc = reg_o; o6_X = reg_o; Enable sign a; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_38 =>
            -- reg_a = a4_X; reg_b = a3_X; reg_acc = reg_o >> 272; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "111";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_39 =>
            -- reg_a = a5_X; reg_b = a2_X; reg_acc = reg_o; o7_X = reg_o; Enable sign a; operation : 2*a*b + acc; Increase base address o;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "111";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '1';
        when square_direct_40 =>
            -- reg_a = a4_X; reg_b = a4_X; reg_acc = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_41 =>
            -- reg_a = a5_X; reg_b = a3_X; reg_acc = reg_o; o8_X = reg_o; Enable sign a; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_42 =>
            -- reg_a = a5_X; reg_b = a4_X; reg_acc = reg_o >> 272; o9_X = reg_o; Enable sign a; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_43 =>
            -- reg_a = a5_X; reg_b = a5_X; reg_acc = reg_o >> 272; o10_X = reg_o; o11_X = reg_o >> 272; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_45 =>
            -- -- Other cases
            -- reg_a = a5_X; reg_b = a0_X; reg_acc = reg_o; o5_X = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_46 =>
            -- reg_a = a3_X; reg_b = a3_X; reg_acc = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_47 =>
            -- reg_a = a4_X; reg_b = a2_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_48 =>
            -- reg_a = a5_X; reg_b = a1_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_49 =>
            -- -- In case of size 7
            -- reg_a = a6_X; reg_b = a0_X; reg_acc = reg_o; o6_X = reg_o; Enable sign a; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_50 =>
            -- reg_a = a4_X; reg_b = a3_X; reg_acc = reg_o >> 272; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "111";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_51 =>
            -- reg_a = a5_X; reg_b = a2_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "111";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_52 =>
            -- reg_a = a6_X; reg_b = a1_X; reg_acc = reg_o; o7_X = reg_o; Enable sign a; operation : 2*a*b + acc; Increase base address o;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "111";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '1';
        when square_direct_53 =>
            -- reg_a = a4_X; reg_b = a4_X; reg_acc = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_54 =>
            -- reg_a = a5_X; reg_b = a3_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_55 =>
            -- reg_a = a6_X; reg_b = a2_X; reg_acc = reg_o; o8_X = reg_o; Enable sign a; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_56 =>
            -- reg_a = a5_X; reg_b = a4_X; reg_acc = reg_o >> 272; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_57 =>
            -- reg_a = a6_X; reg_b = a3_X; reg_acc = reg_o; o9_X = reg_o; Enable sign a; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_58 =>
            -- reg_a = a5_X; reg_b = a5_X; reg_acc = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_59 =>
            -- reg_a = a6_X; reg_b = a4_X; reg_acc = reg_o; o10_X = reg_o; Enable sign a; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_60 =>
            -- reg_a = a6_X; reg_b = a5_X; reg_acc = reg_o >> 272; o11_X = reg_o; Enable sign a; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_61 =>
            -- reg_a = a6_X; reg_b = a6_X; reg_acc = reg_o >> 272; o12_X = reg_o; o13_X = reg_o >> 272; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_63 =>
            -- -- In case of size 8
            -- reg_a = a6_X; reg_b = a0_X; reg_acc = reg_o; o6_X = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_64 =>
            -- reg_a = a4_X; reg_b = a3_X; reg_acc = reg_o >> 272; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "111";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_65 =>
            -- reg_a = a5_X; reg_b = a2_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "111";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_66 =>
            -- reg_a = a6_X; reg_b = a1_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "111";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_67 =>
            -- reg_a = a7_X; reg_b = a0_X; reg_acc = reg_o; o7_X = reg_o; Enable sign a; operation : 2*a*b + acc; Increase base address o;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "111";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '1';
        when square_direct_68 =>
            -- reg_a = a4_X; reg_b = a4_X; reg_acc = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_69 =>
            -- reg_a = a5_X; reg_b = a3_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_70 =>
            -- reg_a = a6_X; reg_b = a2_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_71 =>
            -- reg_a = a7_X; reg_b = a1_X; reg_acc = reg_o; o8_X = reg_o; Enable sign a; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_72 =>
            -- reg_a = a5_X; reg_b = a4_X; reg_acc = reg_o >> 272; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_73 =>
            -- reg_a = a6_X; reg_b = a3_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_74 =>
            -- reg_a = a7_X; reg_b = a2_X; reg_acc = reg_o; o9_X = reg_o; Enable sign a; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_75 =>
            -- reg_a = a5_X; reg_b = a5_X; reg_acc = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_76 =>
            -- reg_a = a6_X; reg_b = a4_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_77 =>
            -- reg_a = a7_X; reg_b = a3_X; reg_acc = reg_o; o10_X = reg_o; Enable sign a; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_78 =>
            -- reg_a = a6_X; reg_b = a5_X; reg_acc = reg_o >> 272; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_79 =>
            -- reg_a = a7_X; reg_b = a4_X; reg_acc = reg_o; o11_X = reg_o; Enable sign a; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_80 =>
            -- reg_a = a6_X; reg_b = a6_X; reg_acc = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_81 =>
            -- reg_a = a7_X; reg_b = a5_X; reg_acc = reg_o; o12_X = reg_o; Enable sign a; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_82 =>
            -- reg_a = a7_X; reg_b = a6_X; reg_acc = reg_o >> 272; o13_X = reg_o; Enable sign a; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_83 =>
            -- reg_a = a7_X; reg_b = a7_X; reg_acc = reg_o >> 272; o14_X = reg_o; o15_X = reg_o >> 272; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
            
            
            
        when multiplication_with_reduction_0 =>
            -- -- In case of size 1
            -- reg_a = a0_X; reg_b = b0_X; reg_acc = 0; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_1 =>
            -- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o0_X = reg_y; operation : keep accumulator;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "11";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "10";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "11";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '1';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_2 =>
            -- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "01";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_3 =>
            -- reg_a = 0; reg_b = 0; reg_acc = reg_o >> 272; o0_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "11";
            next_mac_clear_reg_b <= '1';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_5 =>
            -- -- In case of sizes 2, 3, 4, 5, 6, 7, 8
            -- reg_a = a0_X; reg_b = b0_X; reg_acc = 0; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_6 =>
            -- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o0_X = reg_y; operation : keep accumulator;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "11";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "10";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "11";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '1';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_7 =>
            -- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "01";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_8 =>
            --reg_a = o0_X; reg_b = prime1; reg_acc = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_9 =>
            -- -- In case of size 2
            -- reg_a = a0_X; reg_b = b1_X; reg_acc = reg_o; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_10 =>
            -- reg_a = a1_X; reg_b = b0_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_11 =>
            -- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o1_X = reg_y; operation : keep accumulator;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "11";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "10";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "11";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '1';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_12 =>
            -- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "01";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_13 =>
            -- reg_a = a1_X; reg_b = b1_X; reg_acc = reg_o >> 272; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_14 =>
            -- reg_a = o1_X; reg_b = prime1; reg_acc = reg_o; o0_X = reg_o; o1_X = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_16 =>
            -- -- Other cases
            -- reg_a = a0_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_17 =>
            -- reg_a = a1_X; reg_b = b0_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_18 =>
            -- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o1_X = reg_y; operation : keep accumulator;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "11";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "10";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "11";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '1';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_19 =>
            -- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "01";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_20 =>
            -- reg_a = o0_X; reg_b = prime2; reg_acc = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_21 =>
            -- reg_a = a1_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_22 =>
            -- reg_a = o1_X; reg_b = prime1; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_23 =>
            -- -- In case of size 3
            -- reg_a = a0_X; reg_b = b2_X; reg_acc = reg_o; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_24 =>
            -- reg_a = a2_X; reg_b = b0_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_25 =>
            -- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o2_X = reg_y; operation : keep accumulator;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "11";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "10";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "11";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '1';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_26 =>
            -- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "01";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_27 =>
            -- reg_a = a1_X; reg_b = b2_X; reg_acc = reg_o >> 272; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_28 =>
            -- reg_a = o1_X; reg_b = prime2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_29 =>
            -- reg_a = a2_X; reg_b = b1_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_30 =>
            -- reg_a = o2_X; reg_b = prime1; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_31 =>
            -- reg_a = a2_X; reg_b = b2_X; reg_acc = reg_o >> 272; Enable sign a, b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_32 =>
            -- reg_a = o2_X; reg_b = prime2; reg_acc = reg_o; o1_X = reg_o; o2_X = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_34 =>
            -- -- Other cases
            -- reg_a = a0_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_35 =>
            -- reg_a = a2_X; reg_b = b0_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_36 =>
            -- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o2_X = reg_y; operation : keep accumulator;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "11";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "10";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "11";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '1';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_37 =>
            -- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "01";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_38 =>
            -- reg_a = o0_X; reg_b = prime3; reg_acc = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_39 =>
            -- reg_a = a1_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_40 =>
            -- reg_a = o1_X; reg_b = prime2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_41 =>
            -- reg_a = a2_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_42 =>
            -- reg_a = o2_X; reg_b = prime1; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_43 =>
            -- -- In case of size 4
            -- reg_a = a0_X; reg_b = b3_X; reg_acc = reg_o; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_44 =>
            -- reg_a = a3_X; reg_b = b0_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_45 =>
            -- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o3_X = reg_y; operation : keep accumulator;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "11";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "10";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "11";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '1';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_46 =>
            -- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "01";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_47 =>
            -- reg_a = a1_X; reg_b = b3_X; reg_acc = reg_o >> 272; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_48 =>
            -- reg_a = o1_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_49 =>
            -- reg_a = a2_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_50 =>
            -- reg_a = o2_X; reg_b = prime2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_51 =>
            -- reg_a = a3_X; reg_b = b1_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_52 =>
            -- reg_a = o3_X; reg_b = prime1; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_53 =>
            -- reg_a = a2_X; reg_b = b3_X; reg_acc = reg_o >> 272; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_54 =>
            -- reg_a = o2_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_55 =>
            -- reg_a = a3_X; reg_b = b2_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_56 =>
            -- reg_a = o3_X; reg_b = prime2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_57 =>
            -- reg_a = a3_X; reg_b = b3_X; reg_acc = reg_o >> 272; Enable sign a, b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_58 =>
            -- reg_a = o3_X; reg_b = prime3; reg_acc = reg_o; o2_X = reg_o; o3_0 = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_60 =>
            -- -- Other cases
            -- reg_a = a0_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_61 =>
            -- reg_a = a3_X; reg_b = b0_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_62 =>
            -- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o3_X = reg_y; operation : keep accumulator;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "11";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "10";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "11";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '1';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_63 =>
            -- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "01";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_64 =>
            -- reg_a = o0_X; reg_b = prime4; reg_acc = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_65 =>
            -- reg_a = a1_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_66 =>
            -- reg_a = o1_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_67 =>
            -- reg_a = a2_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_68 =>
            -- reg_a = o2_X; reg_b = prime2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_69 =>
            -- reg_a = a3_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_70 =>
            -- reg_a = o3_X; reg_b = prime1; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_71 =>
            -- -- In case of size 5
            -- reg_a = a0_X; reg_b = b4_X; reg_acc = reg_o; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_72 =>
            -- reg_a = a4_X; reg_b = b0_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_73 =>
            -- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o4_X = reg_y; operation : keep accumulator;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "11";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "10";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "11";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '1';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_74 =>
            -- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "01";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_75 =>
            -- reg_a = a1_X; reg_b = b4_X; reg_acc = reg_o >> 272; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_76 =>
            -- reg_a = o1_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_77 =>
            -- reg_a = a2_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_78 =>
            -- reg_a = o2_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_79 =>
            -- reg_a = a3_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_80 =>
            -- reg_a = o3_X; reg_b = prime2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_81 =>
            -- reg_a = a4_X; reg_b = b1_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_82 =>
            -- reg_a = o4_X; reg_b = prime1; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_83 =>
            -- reg_a = a2_X; reg_b = b4_X; reg_acc = reg_o >> 272; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_84 =>
            -- reg_a = o2_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_85 =>
            -- reg_a = a3_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_86 =>
            -- reg_a = o3_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_87 =>
            -- reg_a = a4_X; reg_b = b2_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_88 =>
            -- reg_a = o4_X; reg_b = prime2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_89 =>
            -- reg_a = a3_X; reg_b = b4_X; reg_acc = reg_o >> 272; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_90 =>
            -- reg_a = o3_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_91 =>
            -- reg_a = a4_X; reg_b = b3_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_92 =>
            -- reg_a = o4_X; reg_b = prime3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_93 =>
            -- reg_a = a4_X; reg_b = b4_X; reg_acc = reg_o >> 272; Enable sign a, b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_94 =>
            -- reg_a = o4_X; reg_b = prime4; reg_acc = reg_o; o3_X = reg_o; o4_0 = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_96 =>
            -- -- Other cases
            -- reg_a = a0_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_97 =>
            -- reg_a = a4_X; reg_b = b0_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_98 =>
            -- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o4_X = reg_y; operation : keep accumulator;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "11";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "10";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "11";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '1';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_99 =>
            -- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "01";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_100 =>
            -- reg_a = o0_X; reg_b = prime5; reg_acc = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_101 =>
            -- reg_a = a1_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_102 =>
            -- reg_a = o1_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_103 =>
            -- reg_a = a2_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_104 =>
            -- reg_a = o2_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_105 =>
            -- reg_a = a3_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_106 =>
            -- reg_a = o3_X; reg_b = prime2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_107 =>
            -- reg_a = a4_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_108 =>
            -- reg_a = o4_X; reg_b = prime1; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_109 =>
            -- -- In case of size 6
            -- reg_a = a0_X; reg_b = b5_X; reg_acc = reg_o; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_110 =>
            -- reg_a = a5_X; reg_b = b0_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_111 =>
            -- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o5_X = reg_y; operation : keep accumulator;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "11";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "10";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "11";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '1';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_112 =>
            -- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "01";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_113 =>
            -- reg_a = a1_X; reg_b = b5_X; reg_acc = reg_o >> 272; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_114 =>
            -- reg_a = o1_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_115 =>
            -- reg_a = a2_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_116 =>
            -- reg_a = o2_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_117 =>
            -- reg_a = a3_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_118 =>
            -- reg_a = o3_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_119 =>
            -- reg_a = a4_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_120 =>
            -- reg_a = o4_X; reg_b = prime2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_121 =>
            -- reg_a = a5_X; reg_b = b1_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_122 =>
            -- reg_a = o5_X; reg_b = prime1; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_123 =>
            -- reg_a = a2_X; reg_b = b5_X; reg_acc = reg_o >> 272; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_124 =>
            -- reg_a = o2_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_125 =>
            -- reg_a = a3_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_126 =>
            -- reg_a = o3_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_127 =>
            -- reg_a = a4_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_128 =>
            -- reg_a = o4_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_129 =>
            -- reg_a = a5_X; reg_b = b2_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_130 =>
            -- reg_a = o5_X; reg_b = prime2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_131 =>
            -- reg_a = a3_X; reg_b = b5_X; reg_acc = reg_o >> 272; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_132 =>
            -- reg_a = o3_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_133 =>
            -- reg_a = a4_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_134 =>
            -- reg_a = o4_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_135 =>
            -- reg_a = a5_X; reg_b = b3_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_136 =>
            -- reg_a = o5_X; reg_b = prime3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_137 =>
            -- reg_a = a4_X; reg_b = b5_X; reg_acc = reg_o >> 272; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_138 =>
            -- reg_a = o4_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_139 =>
            -- reg_a = a5_X; reg_b = b4_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_140 =>
            -- reg_a = o5_X; reg_b = prime4; reg_acc = reg_o; o3_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_141 =>
            -- reg_a = a5_X; reg_b = b5_X; reg_acc = reg_o >> 272; Enable sign a, b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_142 =>
            -- reg_a = o5_X; reg_b = prime5; reg_acc = reg_o; o4_X = reg_o; o5_0 = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_144 =>
            -- -- Other cases
            -- reg_a = a0_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_145 =>
            -- reg_a = a5_X; reg_b = b0_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_146 =>
            -- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o5_X = reg_y; operation : keep accumulator;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "11";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "10";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "11";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '1';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_147 =>
            -- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "01";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_148 =>
            -- reg_a = o0_X; reg_b = prime6; reg_acc = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_149 =>
            -- reg_a = a1_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_150 =>
            -- reg_a = o1_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_151 =>
            -- reg_a = a2_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_152 =>
            -- reg_a = o2_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_153 =>
            -- reg_a = a3_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_154 =>
            -- reg_a = o3_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_155 =>
            -- reg_a = a4_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_156 =>
            -- reg_a = o4_X; reg_b = prime2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_157 =>
            -- reg_a = a5_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_158 =>
            -- reg_a = o5_X; reg_b = prime1; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_159 =>
            -- -- In case of size 7
            -- reg_a = a0_X; reg_b = b6_X; reg_acc = reg_o; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_160 =>
            -- reg_a = a6_X; reg_b = b0_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_161 =>
            -- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o6_X = reg_y; operation : keep accumulator;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "11";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "10";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "11";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '1';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_162 =>
            -- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "01";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_163 =>
            -- reg_a = a1_X; reg_b = b6_X; reg_acc = reg_o >> 272; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_164 =>
            -- reg_a = o1_X; reg_b = prime6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_165 =>
            -- reg_a = a2_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_166 =>
            -- reg_a = o2_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_167 =>
            -- reg_a = a3_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_168 =>
            -- reg_a = o3_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_169 =>
            -- reg_a = a4_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_170 =>
            -- reg_a = o4_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_171 =>
            -- reg_a = a5_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_172 =>
            -- reg_a = o5_X; reg_b = prime2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_173 =>
            -- reg_a = a6_X; reg_b = b1_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_174 =>
            -- reg_a = o6_X; reg_b = prime1; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_175 =>
            -- reg_a = a2_X; reg_b = b6_X; reg_acc = reg_o >> 272; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_176 =>
            -- reg_a = o2_X; reg_b = prime6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_177 =>
            -- reg_a = a3_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_178 =>
            -- reg_a = o3_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_179 =>
            -- reg_a = a4_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_180 =>
            -- reg_a = o4_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_181 =>
            -- reg_a = a5_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_182 =>
            -- reg_a = o5_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_183 =>
            -- reg_a = a6_X; reg_b = b2_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_184 =>
            -- reg_a = o6_X; reg_b = prime2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_185 =>
            -- reg_a = a3_X; reg_b = b6_X; reg_acc = reg_o >> 272; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_186 =>
            -- reg_a = o3_X; reg_b = prime6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_187 =>
            -- reg_a = a4_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_188 =>
            -- reg_a = o4_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_189 =>
            -- reg_a = a5_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_190 =>
            -- reg_a = o5_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_191 =>
            -- reg_a = a6_X; reg_b = b3_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_192 =>
            -- reg_a = o6_X; reg_b = prime3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_193 =>
            -- reg_a = a4_X; reg_b = b6_X; reg_acc = reg_o >> 272; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_194 =>
            -- reg_a = o4_X; reg_b = prime6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_195 =>
            -- reg_a = a5_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_196 =>
            -- reg_a = o5_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_197 =>
            -- reg_a = a6_X; reg_b = b4_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_198 =>
            -- reg_a = o6_X; reg_b = prime4; reg_acc = reg_o; o3_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_199 =>
            -- reg_a = a5_X; reg_b = b6_X; reg_acc = reg_o >> 272; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_200 =>
            -- reg_a = o5_X; reg_b = prime6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_201 =>
            -- reg_a = a6_X; reg_b = b5_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_202 =>
            -- reg_a = o6_X; reg_b = prime5; reg_acc = reg_o; o4_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_203 =>
            -- reg_a = a6_X; reg_b = b6_X; reg_acc = reg_o >> 272; Enable sign a, b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_204 =>
            -- reg_a = o6_X; reg_b = prime6; reg_acc = reg_o; o5_X = reg_o; o6_0 = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_206 =>
            -- -- In case of size 8
            -- reg_a = a0_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_207 =>
            -- reg_a = a6_X; reg_b = b0_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_208 =>
            -- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o6_X = reg_y; operation : keep accumulator;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "11";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "10";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "11";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '1';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_209 =>
            -- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "01";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_210 =>
            -- reg_a = o0_X; reg_b = prime7; reg_acc = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_211 =>
            -- reg_a = a1_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_212 =>
            -- reg_a = o1_X; reg_b = prime6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_213 =>
            -- reg_a = a2_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_214 =>
            -- reg_a = o2_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_215 =>
            -- reg_a = a3_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_216 =>
            -- reg_a = o3_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_217 =>
            -- reg_a = a4_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_218 =>
            -- reg_a = o4_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_219 =>
            -- reg_a = a5_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_220 =>
            -- reg_a = o5_X; reg_b = prime2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_221 =>
            -- reg_a = a6_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_222 =>
            -- reg_a = o6_X; reg_b = prime1; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_223 =>
            -- reg_a = a0_X; reg_b = b7_X; reg_acc = reg_o; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_224 =>
            -- reg_a = a7_X; reg_b = b0_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_225 =>
            -- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o7_X = reg_y; operation : keep accumulator;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "11";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "111";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "10";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "11";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '1';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_226 =>
            -- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "01";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_227 =>
            -- reg_a = a1_X; reg_b = b7_X; reg_acc = reg_o >> 272; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_228 =>
            -- reg_a = o1_X; reg_b = prime7; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_229 =>
            -- reg_a = a2_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_230 =>
            -- reg_a = o2_X; reg_b = prime6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_231 =>
            -- reg_a = a3_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_232 =>
            -- reg_a = o3_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_233 =>
            -- reg_a = a4_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_234 =>
            -- reg_a = o4_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_235 =>
            -- reg_a = a5_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_236 =>
            -- reg_a = o5_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_237 =>
            -- reg_a = a6_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_238 =>
            -- reg_a = o6_X; reg_b = prime2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_239 =>
            -- reg_a = a7_X; reg_b = b1_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_240 =>
            -- reg_a = o7_X; reg_b = prime1; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_241 =>
            -- reg_a = a2_X; reg_b = b7_X; reg_acc = reg_o >> 272; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_242 =>
            -- reg_a = o2_X; reg_b = prime7; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_243 =>
            -- reg_a = a3_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_244 =>
            -- reg_a = o3_X; reg_b = prime6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_245 =>
            -- reg_a = a4_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_246 =>
            -- reg_a = o4_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_247 =>
            -- reg_a = a5_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_248 =>
            -- reg_a = o5_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_249 =>
            -- reg_a = a6_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_250 =>
            -- reg_a = o6_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_251 =>
            -- reg_a = a7_X; reg_b = b2_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_252 =>
            -- reg_a = o7_X; reg_b = prime2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_253 =>
            -- reg_a = a3_X; reg_b = b7_X; reg_acc = reg_o >> 272; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_254 =>
            -- reg_a = o3_X; reg_b = prime7; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_255 =>
            -- reg_a = a4_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_256 =>
            -- reg_a = o4_X; reg_b = prime6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_257 =>
            -- reg_a = a5_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_258 =>
            -- reg_a = o5_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_259 =>
            -- reg_a = a6_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_260 =>
            -- reg_a = o6_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_261 =>
            -- reg_a = a7_X; reg_b = b3_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_262 =>
            -- reg_a = o7_X; reg_b = prime3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_263 =>
            -- reg_a = a4_X; reg_b = b7_X; reg_acc = reg_o >> 272; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_264 =>
            -- reg_a = o4_X; reg_b = prime7; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_265 =>
            -- reg_a = a5_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_266 =>
            -- reg_a = o5_X; reg_b = prime6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_267 =>
            -- reg_a = a6_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_268 =>
            -- reg_a = o6_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_269 =>
            -- reg_a = a7_X; reg_b = b4_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_270 =>
            -- reg_a = o7_X; reg_b = prime4; reg_acc = reg_o; o3_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_271 =>
            -- reg_a = a5_X; reg_b = b7_X; reg_acc = reg_o >> 272; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_272 =>
            -- reg_a = o5_X; reg_b = prime7; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_273 =>
            -- reg_a = a6_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_274 =>
            -- reg_a = o6_X; reg_b = prime6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_275 =>
            -- reg_a = a7_X; reg_b = b5_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_276 =>
            -- reg_a = o7_X; reg_b = prime5; reg_acc = reg_o; o4_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_277 =>
            -- reg_a = a6_X; reg_b = b7_X; reg_acc = reg_o >> 272; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_278 =>
            -- reg_a = o6_X; reg_b = prime7; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_279 =>
            -- reg_a = a7_X; reg_b = b6_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_280 =>
            -- reg_a = o7_X; reg_b = prime6; reg_acc = reg_o; o5_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_281 =>
            -- reg_a = a7_X; reg_b = b7_X; reg_acc = reg_o >> 272; Enable sign a, b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_282 =>
            -- reg_a = o7_X; reg_b = prime7; reg_acc = reg_o; o6_X = reg_o; o7_0 = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_0 =>
            -- -- In case of size 1
            -- reg_a = a0_X; reg_b = b0_X; reg_acc = 0; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1 =>
            -- reg_a = 0; reg_b = 0; reg_acc = reg_o >> 272; o0_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "11";
            next_mac_clear_reg_b <= '1';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3 =>
            -- -- In case of sizes 2, 3, 4
            -- reg_a = a0_X; reg_b = b0_X; reg_acc = 0; o0_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_4 =>
            -- -- In case of size 2
            -- reg_a = a0_X; reg_b = b1_X; reg_acc = reg_o >> 272; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_5 =>
            -- reg_a = o0_X; reg_b = primeSP1; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_6 =>
            -- reg_a = a1_X; reg_b = b0_X; reg_acc = reg_o; o1_X = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_7 =>
            -- reg_a = a1_X; reg_b = b1_X; reg_acc = reg_o >> 272; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_8 =>
            -- reg_a = o1_X; reg_b = primeSP1; reg_acc = reg_o; o0_X = reg_o; o1_X = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_10 =>
            -- -- In case of sizes 3, 4
            -- reg_a = a0_X; reg_b = b1_X; reg_acc = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_11 =>
            -- reg_a = o0_X; reg_b = primeSP1; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_12 =>
            -- reg_a = a1_X; reg_b = b0_X; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_13 =>
            -- reg_a = o0_X; reg_b = primeSP2; reg_acc = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_14 =>
            -- reg_a = a1_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_15 =>
            -- reg_a = o1_X; reg_b = primeSP1; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_16 =>
            -- -- In case of size 3
            -- reg_a = a0_X; reg_b = b2_X; reg_acc = reg_o; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_17 =>
            -- reg_a = a2_X; reg_b = b0_X; reg_acc = reg_o; o2_X = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_18 =>
            -- reg_a = a1_X; reg_b = b2_X; reg_acc = reg_o >> 272; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_19 =>
            -- reg_a = o1_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_20 =>
            -- reg_a = a2_X; reg_b = b1_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_21 =>
            -- reg_a = o2_X; reg_b = primeSP1; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_22 =>
            -- reg_a = a2_X; reg_b = b2_X; reg_acc = reg_o >> 272; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_23 =>
            -- reg_a = o2_X; reg_b = primeSP2; reg_acc = reg_o; o1_X = reg_o; o2_X = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_25 =>
            -- -- In case of size 4
            -- reg_a = a0_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_26 =>
            -- reg_a = a2_X; reg_b = b0_X; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_27 =>
            -- reg_a = o0_X; reg_b = primeSP3; reg_acc = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_28 =>
            -- reg_a = a1_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_29 =>
            -- reg_a = o1_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_30 =>
            -- reg_a = a2_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_31 =>
            -- reg_a = o2_X; reg_b = primeSP1; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_32 =>
            -- reg_a = a0_X; reg_b = b3_X; reg_acc = reg_o; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_33 =>
            -- reg_a = a3_X; reg_b = b0_X; reg_acc = reg_o; o3_X = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_34 =>
            -- reg_a = a1_X; reg_b = b3_X; reg_acc = reg_o >> 272; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_35 =>
            -- reg_a = o1_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_36 =>
            -- reg_a = a2_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_37 =>
            -- reg_a = o2_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_38 =>
            -- reg_a = a3_X; reg_b = b1_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_39 =>
            -- reg_a = o3_X; reg_b = primeSP1; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_40 =>
            -- reg_a = a2_X; reg_b = b3_X; reg_acc = reg_o >> 272; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_41 =>
            -- reg_a = o2_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_42 =>
            -- reg_a = a3_X; reg_b = b2_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_43 =>
            -- reg_a = o3_X; reg_b = primeSP2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_44 =>
            -- reg_a = a3_X; reg_b = b3_X; reg_acc = reg_o >> 272; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_45 =>
            -- reg_a = o3_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; o3_X = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_47 =>
            -- -- In case of sizes 5, 6
            -- reg_a = a0_X; reg_b = b0_X; reg_acc = 0; o0_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_48 =>
            -- reg_a = a0_X; reg_b = b1_X; reg_acc = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_49 =>
            -- reg_a = a1_X; reg_b = b0_X; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_50 =>
            -- reg_a = o0_X; reg_b = primeSP2; reg_acc = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_51 =>
            -- reg_a = a1_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_52 =>
            -- reg_a = a0_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_53 =>
            -- reg_a = a2_X; reg_b = b0_X; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_54 =>
            -- reg_a = o0_X; reg_b = primeSP3; reg_acc = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_55 =>
            -- reg_a = a1_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_56 =>
            -- reg_a = o1_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_57 =>
            -- reg_a = a2_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_58 =>
            -- reg_a = a0_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_59 =>
            -- reg_a = a3_X; reg_b = b0_X; reg_acc = reg_o; o3_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_60 =>
            -- reg_a = o0_X; reg_b = primeSP4; reg_acc = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_61 =>
            -- reg_a = a1_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_62 =>
            -- reg_a = o1_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_63 =>
            -- reg_a = a2_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_64 =>
            -- reg_a = o2_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_65 =>
            -- reg_a = a3_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_66 =>
            -- In case of size 5
            -- reg_a = a0_X; reg_b = b4_X; reg_acc = reg_o; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_67 =>
            -- reg_a = a4_X; reg_b = b0_X; reg_acc = reg_o; o4_X = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_68 =>
            -- reg_a = a1_X; reg_b = b4_X; reg_acc = reg_o >> 272; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_69 =>
            -- reg_a = o1_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_70 =>
            -- reg_a = a2_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_71 =>
            -- reg_a = o2_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_72 =>
            -- reg_a = a3_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_73 =>
            -- reg_a = o3_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_74 =>
            -- reg_a = a4_X; reg_b = b1_X; reg_acc = reg_o; o0_X = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_75 =>
            -- reg_a = a2_X; reg_b = b4_X; reg_acc = reg_o >> 272; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_76 =>
            -- reg_a = o2_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_77 =>
            -- reg_a = a3_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_78 =>
            -- reg_a = o3_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_79 =>
            -- reg_a = a4_X; reg_b = b2_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_80 =>
            -- reg_a = o4_X; reg_b = primeSP2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_81 =>
            -- reg_a = a3_X; reg_b = b4_X; reg_acc = reg_o >> 272; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_82 =>
            -- reg_a = o3_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_83 =>
            -- reg_a = a4_X; reg_b = b3_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_84 =>
            -- reg_a = o4_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_85 =>
            -- reg_a = a4_X; reg_b = b4_X; reg_acc = reg_o >> 272; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_86 =>
            -- reg_a = o4_X; reg_b = primeSP4; reg_acc = reg_o; o3_X = reg_o; o4_X = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_88 =>
            -- -- In case of size 6
            -- reg_a = a0_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_89 =>
            -- reg_a = a4_X; reg_b = b0_X; reg_acc = reg_o; o4_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_90 =>
            -- reg_a = o0_X; reg_b = primeSP5; reg_acc = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_91 =>
            -- reg_a = a1_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_92 =>
            -- reg_a = o1_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_93 =>
            -- reg_a = a2_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_94 =>
            -- reg_a = o2_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_95 =>
            -- reg_a = a3_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_96 =>
            -- reg_a = o3_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_97 =>
            -- reg_a = a4_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_98 =>
            -- reg_a = a0_X; reg_b = b5_X; reg_acc = reg_o; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_99 =>
            -- reg_a = a5_X; reg_b = b0_X; reg_acc = reg_o; o5_X = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_100 =>
            -- reg_a = a1_X; reg_b = b5_X; reg_acc = reg_o >> 272; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_101 =>
            -- reg_a = o1_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_102 =>
            -- reg_a = a2_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_103 =>
            -- reg_a = o2_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_104 =>
            -- reg_a = a3_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_105 =>
            -- reg_a = o3_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_106 =>
            -- reg_a = a4_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_107 =>
            -- reg_a = o4_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_108 =>
            -- reg_a = a5_X; reg_b = b1_X; reg_acc = reg_o; o0_X = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_109 =>
            -- reg_a = a2_X; reg_b = b5_X; reg_acc = reg_o >> 272; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_110 =>
            -- reg_a = o2_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_111 =>
            -- reg_a = a3_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_112 =>
            -- reg_a = o3_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_113 =>
            -- reg_a = a4_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_114 =>
            -- reg_a = o4_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_115 =>
            -- reg_a = a5_X; reg_b = b2_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_116 =>
            -- reg_a = o5_X; reg_b = primeSP2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_117 =>
            -- reg_a = a3_X; reg_b = b5_X; reg_acc = reg_o >> 272; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_118 =>
            -- reg_a = o3_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_119 =>
            -- reg_a = a4_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_120 =>
            -- reg_a = o4_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_121 =>
            -- reg_a = a5_X; reg_b = b3_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_122 =>
            -- reg_a = o5_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_123 =>
            -- reg_a = a4_X; reg_b = b5_X; reg_acc = reg_o >> 272; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_124 =>
            -- reg_a = o4_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_125 =>
            -- reg_a = a5_X; reg_b = b4_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_126 =>
            -- reg_a = o5_X; reg_b = primeSP4; reg_acc = reg_o; o3_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_127 =>
            -- reg_a = a5_X; reg_b = b5_X; reg_acc = reg_o >> 272; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_128 =>
            -- reg_a = o5_X; reg_b = primeSP5; reg_acc = reg_o; o4_X = reg_o; o5_X = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_130 =>
            -- -- In case of sizes 7, 8
            -- reg_a = a0_X; reg_b = b0_X; reg_acc = 0; o0_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_131 =>
            -- reg_a = a0_X; reg_b = b1_X; reg_acc = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_132 =>
            -- reg_a = a1_X; reg_b = b0_X; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_133 =>
            -- reg_a = a1_X; reg_b = b1_X; reg_acc = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_134 =>
            -- reg_a = a0_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_135 =>
            -- reg_a = a2_X; reg_b = b0_X; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_136 =>
            -- reg_a = o0_X; reg_b = primeSP3; reg_acc = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_137 =>
            -- reg_a = a1_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_138 =>
            -- reg_a = a2_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_139 =>
            -- reg_a = a0_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_140 =>
            -- reg_a = a3_X; reg_b = b0_X; reg_acc = reg_o; o3_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_141 =>
            -- reg_a = o0_X; reg_b = primeSP4; reg_acc = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_142 =>
            -- reg_a = a1_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_143 =>
            -- reg_a = o1_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_144 =>
            -- reg_a = a2_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_145 =>
            -- reg_a = a3_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_146 =>
            -- reg_a = a0_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_147 =>
            -- reg_a = a4_X; reg_b = b0_X; reg_acc = reg_o; o4_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_148 =>
            -- reg_a = o0_X; reg_b = primeSP5; reg_acc = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_149 =>
            -- reg_a = a1_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_150 =>
            -- reg_a = o1_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_151 =>
            -- reg_a = a2_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_152 =>
            -- reg_a = o2_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_153 =>
            -- reg_a = a3_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_154 =>
            -- reg_a = a4_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_155 =>
            -- reg_a = a0_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_156 =>
            -- reg_a = a5_X; reg_b = b0_X; reg_acc = reg_o; o5_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_157 =>
            -- reg_a = o0_X; reg_b = primeSP6; reg_acc = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_158 =>
            -- reg_a = a1_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_159 =>
            -- reg_a = o1_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_160 =>
            -- reg_a = a2_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_161 =>
            -- reg_a = o2_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_162 =>
            -- reg_a = a3_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_163 =>
            -- reg_a = o3_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_164 =>
            -- reg_a = a4_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_165 =>
            -- reg_a = a5_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_166 =>
            -- -- In case of size 7
            -- reg_a = a0_X; reg_b = b6_X; reg_acc = reg_o; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_167 =>
            -- reg_a = a6_X; reg_b = b0_X; reg_acc = reg_o; o6_X = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_168 =>
            -- reg_a = a1_X; reg_b = b6_X; reg_acc = reg_o >> 272; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_169 =>
            -- reg_a = o1_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_170 =>
            -- reg_a = a2_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_171 =>
            -- reg_a = o2_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_172 =>
            -- reg_a = a3_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_173 =>
            -- reg_a = o3_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_174 =>
            -- reg_a = a4_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_175 =>
            -- reg_a = o4_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_176 =>
            -- reg_a = a5_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_177 =>
            -- reg_a = a6_X; reg_b = b1_X; reg_acc = reg_o; o0_X = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_178 =>
            -- reg_a = a2_X; reg_b = b6_X; reg_acc = reg_o >> 272; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_179 =>
            -- reg_a = o2_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_180 =>
            -- reg_a = a3_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_181 =>
            -- reg_a = o3_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_182 =>
            -- reg_a = a4_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_183 =>
            -- reg_a = o4_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_184 =>
            -- reg_a = a5_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_185 =>
            -- reg_a = o5_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_186 =>
            -- reg_a = a6_X; reg_b = b2_X; reg_acc = reg_o; o1_X = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_187 =>
            -- reg_a = a3_X; reg_b = b6_X; reg_acc = reg_o >> 272; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_188 =>
            -- reg_a = o3_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_189 =>
            -- reg_a = a4_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_190 =>
            -- reg_a = o4_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_191 =>
            -- reg_a = a5_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_192 =>
            -- reg_a = o5_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_193 =>
            -- reg_a = a6_X; reg_b = b3_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_194 =>
            -- reg_a = o6_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_195 =>
            -- reg_a = a4_X; reg_b = b6_X; reg_acc = reg_o >> 272; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_196 =>
            -- reg_a = o4_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_197 =>
            -- reg_a = a5_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_198 =>
            -- reg_a = o5_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_199 =>
            -- reg_a = a6_X; reg_b = b4_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_200 =>
            -- reg_a = o6_X; reg_b = primeSP4; reg_acc = reg_o; o3_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_201 =>
            -- reg_a = a5_X; reg_b = b6_X; reg_acc = reg_o >> 272; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_202 =>
            -- reg_a = o5_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_203 =>
            -- reg_a = a6_X; reg_b = b5_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_204 =>
            -- reg_a = o6_X; reg_b = primeSP5; reg_acc = reg_o; o4_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_205 =>
            -- reg_a = a6_X; reg_b = b6_X; reg_acc = reg_o >> 272; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_206 =>
            -- reg_a = o6_X; reg_b = primeSP6; reg_acc = reg_o; o5_X = reg_o; o6_X = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_208 =>
            -- -- In case of size 8
            -- reg_a = a0_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_209 =>
            -- reg_a = a6_X; reg_b = b0_X; reg_acc = reg_o; o6_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_210 =>
            -- reg_a = o0_X; reg_b = primeSP7; reg_acc = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_211 =>
            -- reg_a = a1_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_212 =>
            -- reg_a = o1_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_213 =>
            -- reg_a = a2_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_214 =>
            -- reg_a = o2_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_215 =>
            -- reg_a = a3_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_216 =>
            -- reg_a = o3_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_217 =>
            -- reg_a = a4_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_218 =>
            -- reg_a = o4_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_219 =>
            -- reg_a = a5_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_220 =>
            -- reg_a = a6_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_221 =>
            -- reg_a = a0_X; reg_b = b7_X; reg_acc = reg_o; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_222 =>
            -- reg_a = a7_X; reg_b = b0_X; reg_acc = reg_o; o7_X = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "111";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_223 =>
            -- reg_a = a1_X; reg_b = b7_X; reg_acc = reg_o >> 272; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_224 =>
            -- reg_a = o1_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_225 =>
            -- reg_a = a2_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_226 =>
            -- reg_a = o2_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_227 =>
            -- reg_a = a3_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_228 =>
            -- reg_a = o3_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_229 =>
            -- reg_a = a4_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_230 =>
            -- reg_a = o4_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_231 =>
            -- reg_a = a5_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_232 =>
            -- reg_a = o5_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_233 =>
            -- reg_a = a6_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_234 =>
            -- reg_a = a7_X; reg_b = b1_X; reg_acc = reg_o; o0_X = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_235 =>
            -- reg_a = a2_X; reg_b = b7_X; reg_acc = reg_o >> 272; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_236 =>
            -- reg_a = o2_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_237 =>
            -- reg_a = a3_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_238 =>
            -- reg_a = o3_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_239 =>
            -- reg_a = a4_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_240 =>
            -- reg_a = o4_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_241 =>
            -- reg_a = a5_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_242 =>
            -- reg_a = o5_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_243 =>
            -- reg_a = a6_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_244 =>
            -- reg_a = o6_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_245 =>
            -- reg_a = a7_X; reg_b = b2_X; reg_acc = reg_o; o1_X = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_246 =>
            -- reg_a = a3_X; reg_b = b7_X; reg_acc = reg_o >> 272; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_247 =>
            -- reg_a = o3_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_248 =>
            -- reg_a = a4_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_249 =>
            -- reg_a = o4_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_250 =>
            -- reg_a = a5_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_251 =>
            -- reg_a = o5_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_252 =>
            -- reg_a = a6_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_253 =>
            -- reg_a = o6_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_254 =>
            -- reg_a = a7_X; reg_b = b3_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_255 =>
            -- reg_a = o7_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_256 =>
            -- reg_a = a4_X; reg_b = b7_X; reg_acc = reg_o >> 272; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_257 =>
            -- reg_a = o4_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_258 =>
            -- reg_a = a5_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_259 =>
            -- reg_a = o5_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_260 =>
            -- reg_a = a6_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_261 =>
            -- reg_a = o6_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_262 =>
            -- reg_a = a7_X; reg_b = b4_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_263 =>
            -- reg_a = o7_X; reg_b = primeSP4; reg_acc = reg_o; o3_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_264 =>
            -- reg_a = a5_X; reg_b = b7_X; reg_acc = reg_o >> 272; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_265 =>
            -- reg_a = o5_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_266 =>
            -- reg_a = a6_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_267 =>
            -- reg_a = o6_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_268 =>
            -- reg_a = a7_X; reg_b = b5_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_269 =>
            -- reg_a = o7_X; reg_b = primeSP5; reg_acc = reg_o; o4_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_270 =>
            -- reg_a = a6_X; reg_b = b7_X; reg_acc = reg_o >> 272; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_271 =>
            -- reg_a = o6_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_272 =>
            -- reg_a = a7_X; reg_b = b6_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_273 =>
            -- reg_a = o7_X; reg_b = primeSP6; reg_acc = reg_o; o5_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_274 =>
            -- reg_a = a7_X; reg_b = b7_X; reg_acc = reg_o >> 272; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_275 =>
            -- reg_a = o7_X; reg_b = primeSP7; reg_acc = reg_o; o6_X = reg_o; o7_X = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_0 =>
            -- -- In case of size 1
            -- reg_a = a0_X; reg_b = a0_X; reg_acc = 0; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_1 =>
            -- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o0_X = reg_y; operation : keep accumulator;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "11";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "10";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "11";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '1';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_2 =>
            -- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "01";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_3 =>
            -- reg_a = 0; reg_b = 0; reg_acc = reg_o >> 272; o0_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "11";
            next_mac_clear_reg_b <= '1';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_5 =>
            -- -- In case of 2, 3, 4, 5, 6, 7, 8
            -- reg_a = a0_X; reg_b = a0_X; reg_acc = 0; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_6 =>
            -- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o0_X = reg_y; operation : keep accumulator;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "11";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "10";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "11";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '1';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_7 =>
            -- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "01";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_8 =>
            -- reg_a = o0_X; reg_b = prime1; reg_acc = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_9 =>
            -- -- In case of size 2
            -- reg_a = a0_X; reg_b = a1_X; reg_acc = reg_o; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_10 =>
            -- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o1_X = reg_y; operation : keep accumulator;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "11";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "10";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "11";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '1';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_11 =>
            -- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "01";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_12 =>
            -- reg_a = a1_X; reg_b = a1_X; reg_acc = reg_o >> 272; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_13 =>
            -- reg_a = o1_X; reg_b = prime1; reg_acc = reg_o; o0_X = reg_o; o1_X = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_15 =>
            -- -- Others cases
            -- reg_a = a0_X; reg_b = a1_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_16 =>
            -- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o1_X = reg_y; operation : keep accumulator;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "11";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "10";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "11";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '1';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_17 =>
            -- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "01";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_18 =>
            -- reg_a = o0_X; reg_b = prime2; reg_acc = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_19 =>
            -- reg_a = a1_X; reg_b = a1_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_20 =>
            -- reg_a = o1_X; reg_b = prime1; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_21 =>
            -- -- In case of size 3
            -- reg_a = a0_X; reg_b = a2_X; reg_acc = reg_o; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_22 =>
            -- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o2_X = reg_y; operation : keep accumulator;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "11";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "10";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "11";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '1';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_23 =>
            -- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "01";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_24 =>
            -- reg_a = a1_X; reg_b = a2_X; reg_acc = reg_o >> 272; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_25 =>
            -- reg_a = o1_X; reg_b = prime2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_26 =>
            -- reg_a = o2_X; reg_b = prime1; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_27 =>
            -- reg_a = a2_X; reg_b = a2_X; reg_acc = reg_o >> 272; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_28 =>
            -- reg_a = o2_X; reg_b = prime2; reg_acc = reg_o; o1_X = reg_o; o2_X = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_30 =>
            -- -- Other cases
            -- reg_a = a0_X; reg_b = a2_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_31 =>
            -- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o2_X = reg_y; operation : keep accumulator;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "11";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "10";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "11";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '1';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_32 =>
            -- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "01";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_33 =>
            -- reg_a = o0_X; reg_b = prime3; reg_acc = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_34 =>
            -- reg_a = a1_X; reg_b = a2_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_35 =>
            -- reg_a = o1_X; reg_b = prime2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_36 =>
            -- reg_a = o2_X; reg_b = prime1; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_37 =>
            -- In case of size 4
            -- reg_a = a0_X; reg_b = a3_X; reg_acc = reg_o; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_38 =>
            -- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o3_X = reg_y; operation : keep accumulator;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "11";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "10";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "11";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '1';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_39 =>
            -- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "01";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_40 =>
            -- reg_a = a1_X; reg_b = a3_X; reg_acc = reg_o >> 272; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_41 =>
            -- reg_a = o1_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_42 =>
            -- reg_a = a2_X; reg_b = a2_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_43 =>
            -- reg_a = o2_X; reg_b = prime2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_44 =>
            -- reg_a = o3_X; reg_b = prime1; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_45 =>
            -- reg_a = a2_X; reg_b = a3_X; reg_acc = reg_o >> 272; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_46 =>
            -- reg_a = o2_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_47 =>
            -- reg_a = o3_X; reg_b = prime2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_48 =>
            -- reg_a = a3_X; reg_b = a3_X; reg_acc = reg_o >> 272; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_49 =>
            -- reg_a = o3_X; reg_b = prime3; reg_acc = reg_o; o2_X = reg_o; o3_X = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_51 =>
            -- -- Other cases
            -- reg_a = a0_X; reg_b = a3_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_52 =>
            -- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o3_X = reg_y; operation : keep accumulator;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "11";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "10";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "11";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '1';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_53 =>
            -- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "01";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_54 =>
            -- reg_a = o0_X; reg_b = prime4; reg_acc = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_55 =>
            -- reg_a = a1_X; reg_b = a3_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_56 =>
            -- reg_a = o1_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_57 =>
            -- reg_a = a2_X; reg_b = a2_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_58 =>
            -- reg_a = o2_X; reg_b = prime2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_59 =>
            -- reg_a = o3_X; reg_b = prime1; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_60 =>
            -- -- In case of size 5
            -- reg_a = a0_X; reg_b = a4_X; reg_acc = reg_o; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_61 =>
            -- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o4_X = reg_y; operation : keep accumulator;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "11";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "10";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "11";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '1';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_62 =>
            -- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "01";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_63 =>
            -- reg_a = a1_X; reg_b = a4_X; reg_acc = reg_o >> 272; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_64 =>
            -- reg_a = o1_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_65 =>
            -- reg_a = a2_X; reg_b = a3_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_66 =>
            -- reg_a = o2_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_67 =>
            -- reg_a = o3_X; reg_b = prime2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_68 =>
            -- reg_a = o4_X; reg_b = prime1; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_69 =>
            -- reg_a = a2_X; reg_b = a4_X; reg_acc = reg_o >> 272; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_70 =>
            -- reg_a = o2_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_71 =>
            -- reg_a = a3_X; reg_b = a3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_72 =>
            -- reg_a = o3_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_73 =>
            -- reg_a = o4_X; reg_b = prime2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_74 =>
            -- reg_a = a3_X; reg_b = a4_X; reg_acc = reg_o >> 272; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_75 =>
            -- reg_a = o3_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_76 =>
            -- reg_a = o4_X; reg_b = prime3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_77 =>
            -- reg_a = a4_X; reg_b = a4_X; reg_acc = reg_o >> 272; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_78 =>
            -- reg_a = o4_X; reg_b = prime4; reg_acc = reg_o; o3_X = reg_o; o4_X = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_80 =>
            -- -- Other cases
            -- reg_a = a0_X; reg_b = a4_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_81 =>
            -- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o4_X = reg_y; operation : keep accumulator;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "11";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "10";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "11";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '1';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_82 =>
            -- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "01";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_83 =>
            -- reg_a = o0_X; reg_b = prime5; reg_acc = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_84 =>
            -- reg_a = a1_X; reg_b = a4_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_85 =>
            -- reg_a = o1_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_86 =>
            -- reg_a = a2_X; reg_b = a3_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_87 =>
            -- reg_a = o2_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_88 =>
            -- reg_a = o3_X; reg_b = prime2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_89 =>
            -- reg_a = o4_X; reg_b = prime1; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_90 =>
            -- -- In case of size 6
            -- reg_a = a0_X; reg_b = a5_X; reg_acc = reg_o; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_91 =>
            -- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o5_X = reg_y; operation : keep accumulator;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "11";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "10";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "11";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '1';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_92 =>
            -- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "01";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_93 =>
            -- reg_a = a1_X; reg_b = a5_X; reg_acc = reg_o >> 272; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_94 =>
            -- reg_a = o1_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_95 =>
            -- reg_a = a2_X; reg_b = a4_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_96 =>
            -- reg_a = o2_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_97 =>
            -- reg_a = a3_X; reg_b = a3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_98 =>
            -- reg_a = o3_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_99 =>
            -- reg_a = o4_X; reg_b = prime2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_100 =>
            -- reg_a = o5_X; reg_b = prime1; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_101 =>
            -- reg_a = a2_X; reg_b = a5_X; reg_acc = reg_o >> 272; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_102 =>
            -- reg_a = o2_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_103 =>
            -- reg_a = a3_X; reg_b = a4_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_104 =>
            -- reg_a = o3_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_105 =>
            -- reg_a = o4_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_106 =>
            -- reg_a = o5_X; reg_b = prime2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_107 =>
            -- reg_a = a3_X; reg_b = a5_X; reg_acc = reg_o >> 272; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_108 =>
            -- reg_a = o3_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_109 =>
            -- reg_a = a4_X; reg_b = a4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_110 =>
            -- reg_a = o4_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_111 =>
            -- reg_a = o5_X; reg_b = prime3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_112 =>
            -- reg_a = a4_X; reg_b = a5_X; reg_acc = reg_o >> 272; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_113 =>
            -- reg_a = o4_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_114 =>
            -- reg_a = o5_X; reg_b = prime4; reg_acc = reg_o; o3_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_115 =>
            -- reg_a = a5_X; reg_b = a5_X; reg_acc = reg_o >> 272; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_116 =>
            -- reg_a = o5_X; reg_b = prime5; reg_acc = reg_o; o4_X = reg_o; o5_X = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_118 =>
            -- -- Other cases
            -- reg_a = a0_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_119 =>
            -- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o5_X = reg_y; operation : keep accumulator;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "11";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "10";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "11";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '1';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_120 =>
            -- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "01";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_121 =>
            -- reg_a = o0_X; reg_b = prime6; reg_acc = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_122 =>
            -- reg_a = a1_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_123 =>
            -- reg_a = o1_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_124 =>
            -- reg_a = a2_X; reg_b = a4_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_125 =>
            -- reg_a = o2_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_126 =>
            -- reg_a = a3_X; reg_b = a3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_127 =>
            -- reg_a = o3_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_128 =>
            -- reg_a = o4_X; reg_b = prime2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_129 =>
            -- reg_a = o5_X; reg_b = prime1; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_130 =>
            -- -- In case of size 7
            -- reg_a = a0_X; reg_b = a6_X; reg_acc = reg_o; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_131 =>
            -- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o6_X = reg_y; operation : keep accumulator;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "11";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "10";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "11";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '1';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_132 =>
            -- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "01";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_133 =>
            -- reg_a = a1_X; reg_b = a6_X; reg_acc = reg_o >> 272; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_134 =>
            -- reg_a = o1_X; reg_b = prime6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_135 =>
            -- reg_a = a2_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_136 =>
            -- reg_a = o2_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_137 =>
            -- reg_a = a3_X; reg_b = a4_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_138 =>
            -- reg_a = o3_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_139 =>
            -- reg_a = o4_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_140 =>
            -- reg_a = o5_X; reg_b = prime2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_141 =>
            -- reg_a = o6_X; reg_b = prime1; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_142 =>
            -- reg_a = a2_X; reg_b = a6_X; reg_acc = reg_o >> 272; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_143 =>
            -- reg_a = o2_X; reg_b = prime6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_144 =>
            -- reg_a = a3_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_145 =>
            -- reg_a = o3_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_146 =>
            -- reg_a = a4_X; reg_b = a4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_147 =>
            -- reg_a = o4_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_148 =>
            -- reg_a = o5_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_149 =>
            -- reg_a = o6_X; reg_b = prime2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_150 =>
            -- reg_a = a3_X; reg_b = a6_X; reg_acc = reg_o >> 272; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_151 =>
            -- reg_a = o3_X; reg_b = prime6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_152 =>
            -- reg_a = a4_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_153 =>
            -- reg_a = o4_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_154 =>
            -- reg_a = o5_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_155 =>
            -- reg_a = o6_X; reg_b = prime3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_156 =>
            -- reg_a = a4_X; reg_b = a6_X; reg_acc = reg_o >> 272; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_157 =>
            -- reg_a = o4_X; reg_b = prime6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_158 =>
            -- reg_a = a5_X; reg_b = a5_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_159 =>
            -- reg_a = o5_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_160 =>
            -- reg_a = o6_X; reg_b = prime4; reg_acc = reg_o; o3_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_161 =>
            -- reg_a = a5_X; reg_b = a6_X; reg_acc = reg_o >> 272; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_162 =>
            -- reg_a = o5_X; reg_b = prime6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_163 =>
            -- reg_a = o6_X; reg_b = prime5; reg_acc = reg_o; o4_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_164 =>
            -- reg_a = a6_X; reg_b = a6_X; reg_acc = reg_o >> 272; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_165 =>
            -- reg_a = o6_X; reg_b = prime6; reg_acc = reg_o; o5_X = reg_o; o6_X = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_167 =>
            -- -- In case of size 8
            -- reg_a = a0_X; reg_b = a6_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_168 =>
            -- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o6_X = reg_y; operation : keep accumulator;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "11";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "10";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "11";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '1';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_169 =>
            -- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "01";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_170 =>
            -- reg_a = o0_X; reg_b = prime7; reg_acc = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_171 =>
            -- reg_a = a1_X; reg_b = a6_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_172 =>
            -- reg_a = o1_X; reg_b = prime6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_173 =>
            -- reg_a = a2_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_174 =>
            -- reg_a = o2_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_175 =>
            -- reg_a = a3_X; reg_b = a4_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_176 =>
            -- reg_a = o3_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_177 =>
            -- reg_a = o4_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_178 =>
            -- reg_a = o5_X; reg_b = prime2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_179 =>
            -- reg_a = o6_X; reg_b = prime1; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_180 =>
            -- reg_a = a0_X; reg_b = a7_X; reg_acc = reg_o; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_181 =>
            -- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o7_X = reg_y; operation : keep accumulator;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "11";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "111";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "10";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "11";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '1';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_182 =>
            -- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "01";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_183 =>
            -- reg_a = a1_X; reg_b = a7_X; reg_acc = reg_o >> 272; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_184 =>
            -- reg_a = o1_X; reg_b = prime7; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_185 =>
            -- reg_a = a2_X; reg_b = a6_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_186 =>
            -- reg_a = o2_X; reg_b = prime6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_187 =>
            -- reg_a = a3_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_188 =>
            -- reg_a = o3_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_189 =>
            -- reg_a = a4_X; reg_b = a4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_190 =>
            -- reg_a = o4_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_191 =>
            -- reg_a = o5_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_192 =>
            -- reg_a = o6_X; reg_b = prime2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_193 =>
            -- reg_a = o7_X; reg_b = prime1; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_194 =>
            -- reg_a = a2_X; reg_b = a7_X; reg_acc = reg_o >> 272; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_195 =>
            -- reg_a = o2_X; reg_b = prime7; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_196 =>
            -- reg_a = a3_X; reg_b = a6_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_197 =>
            -- reg_a = o3_X; reg_b = prime6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_198 =>
            -- reg_a = a4_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_199 =>
            -- reg_a = o4_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_200 =>
            -- reg_a = o5_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_201 =>
            -- reg_a = o6_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_202 =>
            -- reg_a = o7_X; reg_b = prime2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_203 =>
            -- reg_a = a3_X; reg_b = a7_X; reg_acc = reg_o >> 272; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_204 =>
            -- reg_a = o3_X; reg_b = prime7; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_205 =>
            -- reg_a = a4_X; reg_b = a6_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_206 =>
            -- reg_a = o4_X; reg_b = prime6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_207 =>
            -- reg_a = a5_X; reg_b = a5_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_208 =>
            -- reg_a = o5_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_209 =>
            -- reg_a = o6_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_210 =>
            -- reg_a = o7_X; reg_b = prime3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_211 =>
            -- reg_a = a4_X; reg_b = a7_X; reg_acc = reg_o >> 272; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_212 =>
            -- reg_a = o4_X; reg_b = prime7; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_213 =>
            -- reg_a = a5_X; reg_b = a6_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_214 =>
            -- reg_a = o5_X; reg_b = prime6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_215 =>
            -- reg_a = o6_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_216 =>
            -- reg_a = o7_X; reg_b = prime4; reg_acc = reg_o; o3_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_217 =>
            -- reg_a = a5_X; reg_b = a7_X; reg_acc = reg_o >> 272; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_218 =>
            -- reg_a = o5_X; reg_b = prime7; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_219 =>
            -- reg_a = a6_X; reg_b = a6_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_220 =>
            -- reg_a = o6_X; reg_b = prime6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_221 =>
            -- reg_a = o7_X; reg_b = prime5; reg_acc = reg_o; o4_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_222 =>
            -- reg_a = a6_X; reg_b = a7_X; reg_acc = reg_o >> 272; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_223 =>
            -- reg_a = o6_X; reg_b = prime7; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_224 =>
            -- reg_a = o7_X; reg_b = prime6; reg_acc = reg_o; o5_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_225 =>
            -- reg_a = a7_X; reg_b = a7_X; reg_acc = reg_o >> 272; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_226 =>
            -- reg_a = o7_X; reg_b = prime7; reg_acc = reg_o; o6_X = reg_o; o7_X = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_0 =>
            -- -- In case of size 1
            -- reg_a = a0_X; reg_b = a0_X; reg_acc = 0; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1 =>
            -- reg_a = 0; reg_b = 0; reg_acc = reg_o >> 272; o0_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "11";
            next_mac_clear_reg_b <= '1';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3 =>
            -- -- In case of size 2, 3, 4
            -- reg_a = a0_X; reg_b = a0_X; reg_acc = 0; o0_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_4 =>
            -- reg_a = reg_o; reg_b = primeSP1; reg_acc = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "10";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_5 =>
            -- -- In case of size 2
            -- reg_a = a0_X; reg_b = a1_X; reg_acc = reg_o; o1_X = reg_o; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_6 =>
            -- reg_a = a1_X; reg_b = a1_X; reg_acc = reg_o >> 272; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_7 =>
            -- reg_a = o1_X; reg_b = primeSP1; reg_acc = reg_o; o0_X = reg_o; o1_X = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_9 =>
            -- -- In case of size 3, 4
            -- reg_a = a0_X; reg_b = a1_X; reg_acc = reg_o; o1_X = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_10 =>
            -- reg_a = o0_X; reg_b = primeSP2; reg_acc = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_11 =>
            -- reg_a = a1_X; reg_b = a1_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_12 =>
            -- reg_a = o1_X; reg_b = primeSP1; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_13 =>
            -- -- In case of size 3
            -- reg_a = a0_X; reg_b = a2_X; reg_acc = reg_o; o2_X = reg_o; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_14 =>
            -- reg_a = a1_X; reg_b = a2_X; reg_acc = reg_o >> 272; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_15 =>
            -- reg_a = o1_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_16 =>
            -- reg_a = o2_X; reg_b = primeSP1; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_17 =>
            -- reg_a = a2_X; reg_b = a2_X; reg_acc = reg_o >> 272; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_18 =>
            -- reg_a = o2_X; reg_b = primeSP2; reg_acc = reg_o; o1_X = reg_o; o2_X = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_20 =>
            -- -- In case of size 4
            -- reg_a = a0_X; reg_b = a2_X; reg_acc = reg_o; o2_X = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_21 =>
            -- reg_a = o0_X; reg_b = primeSP3; reg_acc = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_22 =>
            -- reg_a = a1_X; reg_b = a2_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_23 =>
            -- reg_a = o1_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_24 =>
            -- reg_a = o2_X; reg_b = primeSP1; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_25 =>
            -- reg_a = a0_X; reg_b = a3_X; reg_acc = reg_o; o3_X = reg_o; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_26 =>
            -- reg_a = a1_X; reg_b = a3_X; reg_acc = reg_o >> 272; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_27 =>
            -- reg_a = o1_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_28 =>
            -- reg_a = a2_X; reg_b = a2_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_29 =>
            -- reg_a = o2_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_30 =>
            -- reg_a = o3_X; reg_b = primeSP1; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_31 =>
            -- reg_a = a2_X; reg_b = a3_X; reg_acc = reg_o >> 272; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_32 =>
            -- reg_a = o2_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_33 =>
            -- reg_a = o3_X; reg_b = primeSP2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_34 =>
            -- reg_a = a3_X; reg_b = a3_X; reg_acc = reg_o >> 272; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_35 =>
            -- reg_a = o3_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; o3_X = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_37 =>
            -- -- In case of size 5, 6
            -- reg_a = a0_X; reg_b = a0_X; reg_acc = 0; o0_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_38 =>
            -- reg_a = a0_X; reg_b = a1_X; reg_acc = reg_o >> 272; o1_X = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_39 =>
            -- reg_a = o0_X; reg_b = primeSP2; reg_acc = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_40 =>
            -- reg_a = a1_X; reg_b = a1_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_41 =>
            -- reg_a = a0_X; reg_b = a2_X; reg_acc = reg_o; o2_X = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_42 =>
            -- reg_a = o0_X; reg_b = primeSP3; reg_acc = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_43 =>
            -- reg_a = a1_X; reg_b = a2_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_44 =>
            -- reg_a = o1_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_45 =>
            -- reg_a = a0_X; reg_b = a3_X; reg_acc = reg_o; o3_X = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_46 =>
            -- reg_a = o0_X; reg_b = primeSP4; reg_acc = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_47 =>
            -- reg_a = a1_X; reg_b = a3_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_48 =>
            -- reg_a = o1_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_49 =>
            -- reg_a = a2_X; reg_b = a2_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_50 =>
            -- reg_a = o2_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_51 =>
            -- -- In case of size 5
            -- reg_a = a0_X; reg_b = a4_X; reg_acc = reg_o; o4_X = reg_o; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_52 =>
            -- reg_a = a1_X; reg_b = a4_X; reg_acc = reg_o >> 272; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_53 =>
            -- reg_a = o1_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_54 =>
            -- reg_a = a2_X; reg_b = a3_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_55 =>
            -- reg_a = o2_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_56 =>
            -- reg_a = o3_X; reg_b = primeSP2; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_57 =>
            -- reg_a = a2_X; reg_b = a4_X; reg_acc = reg_o >> 272; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_58 =>
            -- reg_a = o2_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_59 =>
            -- reg_a = a3_X; reg_b = a3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_60 =>
            -- reg_a = o3_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_61 =>
            -- reg_a = o4_X; reg_b = primeSP2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_62 =>
            -- reg_a = a3_X; reg_b = a4_X; reg_acc = reg_o >> 272; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_63 =>
            -- reg_a = o3_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_64 =>
            -- reg_a = o4_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_65 =>
            -- reg_a = a4_X; reg_b = a4_X; reg_acc = reg_o >> 272; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_66 =>
            -- reg_a = o4_X; reg_b = primeSP4; reg_acc = reg_o; o3_X = reg_o; o4_X = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_68 =>
            -- -- In case of size 6
            -- reg_a = a0_X; reg_b = a4_X; reg_acc = reg_o; o4_X = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_69 =>
            -- reg_a = o0_X; reg_b = primeSP5; reg_acc = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_70 =>
            -- reg_a = a1_X; reg_b = a4_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_71 =>
            -- reg_a = o1_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_72 =>
            -- reg_a = a2_X; reg_b = a3_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_73 =>
            -- reg_a = o2_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_74 =>
            -- reg_a = o3_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_75 =>
            -- reg_a = a0_X; reg_b = a5_X; reg_acc = reg_o; o5_X = reg_o; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_76 =>
            -- reg_a = a1_X; reg_b = a5_X; reg_acc = reg_o >> 272; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_77 =>
            -- reg_a = o1_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_78 =>
            -- reg_a = a2_X; reg_b = a4_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_79 =>
            -- reg_a = o2_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_80 =>
            -- reg_a = a3_X; reg_b = a3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_81 =>
            -- reg_a = o3_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_82 =>
            -- reg_a = o4_X; reg_b = primeSP2; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_83 =>
            -- reg_a = a2_X; reg_b = a5_X; reg_acc = reg_o >> 272; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_84 =>
            -- reg_a = o2_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_85 =>
            -- reg_a = a3_X; reg_b = a4_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_86 =>
            -- reg_a = o3_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_87 =>
            -- reg_a = o4_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_88 =>
            -- reg_a = o5_X; reg_b = primeSP2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_89 =>
            -- reg_a = a3_X; reg_b = a5_X; reg_acc = reg_o >> 272; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_90 =>
            -- reg_a = o3_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_91 =>
            -- reg_a = a4_X; reg_b = a4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_92 =>
            -- reg_a = o4_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_93 =>
            -- reg_a = o5_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_94 =>
            -- reg_a = a4_X; reg_b = a5_X; reg_acc = reg_o >> 272; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_95 =>
            -- reg_a = o4_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_96 =>
            -- reg_a = o5_X; reg_b = primeSP4; reg_acc = reg_o; o3_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_97 =>
            -- reg_a = a5_X; reg_b = a5_X; reg_acc = reg_o >> 272; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_98 =>
            -- reg_a = o5_X; reg_b = primeSP5; reg_acc = reg_o; o4_X = reg_o; o5_X = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_100 =>
            -- -- In case of size 7, 8
            -- reg_a = a0_X; reg_b = a0_X; reg_acc = 0; o0_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_101 =>
            -- reg_a = a0_X; reg_b = a1_X; reg_acc = reg_o >> 272; o1_X = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_102 =>
            -- reg_a = a1_X; reg_b = a1_X; reg_acc = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_103 =>
            -- reg_a = a0_X; reg_b = a2_X; reg_acc = reg_o; o2_X = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_104 =>
            -- reg_a = o0_X; reg_b = primeSP3; reg_acc = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_105 =>
            -- reg_a = a1_X; reg_b = a2_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_106 =>
            -- reg_a = a0_X; reg_b = a3_X; reg_acc = reg_o; o3_X = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_107 =>
            -- reg_a = o0_X; reg_b = primeSP4; reg_acc = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_108 =>
            -- reg_a = a1_X; reg_b = a3_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_109 =>
            -- reg_a = o1_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_110 =>
            -- reg_a = a2_X; reg_b = a2_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_111 =>
            -- reg_a = a0_X; reg_b = a4_X; reg_acc = reg_o; o4_X = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_112 =>
            -- reg_a = o0_X; reg_b = primeSP5; reg_acc = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_113 =>
            -- reg_a = a1_X; reg_b = a4_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_114 =>
            -- reg_a = o1_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_115 =>
            -- reg_a = a2_X; reg_b = a3_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_116 =>
            -- reg_a = o2_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_117 =>
            -- reg_a = a0_X; reg_b = a5_X; reg_acc = reg_o; o5_X = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_118 =>
            -- reg_a = o0_X; reg_b = primeSP6; reg_acc = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_119 =>
            -- reg_a = a1_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_120 =>
            -- reg_a = o1_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_121 =>
            -- reg_a = a2_X; reg_b = a4_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_122 =>
            -- reg_a = o2_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_123 =>
            -- reg_a = a3_X; reg_b = a3_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_124 =>
            -- reg_a = o3_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_125 =>
            -- -- In case of size 7
            -- reg_a = a0_X; reg_b = a6_X; reg_acc = reg_o; o6_X = reg_o; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_126 =>
            -- reg_a = a1_X; reg_b = a6_X; reg_acc = reg_o >> 272; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_127 =>
            -- reg_a = o1_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_128 =>
            -- reg_a = a2_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_129 =>
            -- reg_a = o2_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_130 =>
            -- reg_a = a3_X; reg_b = a4_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_131 =>
            -- reg_a = o3_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_132 =>
            -- reg_a = o4_X; reg_b = primeSP3; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_133 =>
            -- reg_a = a2_X; reg_b = a6_X; reg_acc = reg_o >> 272; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_134 =>
            -- reg_a = o2_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_135 =>
            -- reg_a = a3_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_136 =>
            -- reg_a = o3_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_137 =>
            -- reg_a = a4_X; reg_b = a4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_138 =>
            -- reg_a = o4_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_139 =>
            -- reg_a = o5_X; reg_b = primeSP3; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_140 =>
            -- reg_a = a3_X; reg_b = a6_X; reg_acc = reg_o >> 272; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_141 =>
            -- reg_a = o3_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_142 =>
            -- reg_a = a4_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_143 =>
            -- reg_a = o4_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_144 =>
            -- reg_a = o5_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_145 =>
            -- reg_a = o6_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_146 =>
            -- reg_a = a4_X; reg_b = a6_X; reg_acc = reg_o >> 272; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_147 =>
            -- reg_a = o4_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_148 =>
            -- reg_a = a5_X; reg_b = a5_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_149 =>
            -- reg_a = o5_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_150 =>
            -- reg_a = o6_X; reg_b = primeSP4; reg_acc = reg_o; o3_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_151 =>
            -- reg_a = a5_X; reg_b = a6_X; reg_acc = reg_o >> 272; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_152 =>
            -- reg_a = o5_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_153 =>
            -- reg_a = o6_X; reg_b = primeSP5; reg_acc = reg_o; o4_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_154 =>
            -- reg_a = a6_X; reg_b = a6_X; reg_acc = reg_o >> 272; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_155 =>
            -- reg_a = o6_X; reg_b = primeSP6; reg_acc = reg_o; o5_X = reg_o; o6_X = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_157 =>
            -- -- In case of size 8
            -- reg_a = a0_X; reg_b = a6_X; reg_acc = reg_o; o6_X = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_158 =>
            -- reg_a = o0_X; reg_b = primeSP7; reg_acc = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_159 =>
            -- reg_a = a1_X; reg_b = a6_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_160 =>
            -- reg_a = o1_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_161 =>
            -- reg_a = a2_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_162 =>
            -- reg_a = o2_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_163 =>
            -- reg_a = a3_X; reg_b = a4_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_164 =>
            -- reg_a = o3_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_165 =>
            -- reg_a = o4_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_166 =>
            -- reg_a = a0_X; reg_b = a7_X; reg_acc = reg_o; o7_X = reg_o; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "111";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_167 =>
            -- reg_a = a1_X; reg_b = a7_X; reg_acc = reg_o >> 272; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_168 =>
            -- reg_a = o1_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_169 =>
            -- reg_a = a2_X; reg_b = a6_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_170 =>
            -- reg_a = o2_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_171 =>
            -- reg_a = a3_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_172 =>
            -- reg_a = o3_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_173 =>
            -- reg_a = a4_X; reg_b = a4_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_174 =>
            -- reg_a = o4_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_175 =>
            -- reg_a = o5_X; reg_b = primeSP3; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_176 =>
            -- reg_a = a2_X; reg_b = a7_X; reg_acc = reg_o >> 272; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_177 =>
            -- reg_a = o2_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_178 =>
            -- reg_a = a3_X; reg_b = a6_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_179 =>
            -- reg_a = o3_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_180 =>
            -- reg_a = a4_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_181 =>
            -- reg_a = o4_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_182 =>
            -- reg_a = o5_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_183 =>
            -- reg_a = o6_X; reg_b = primeSP3; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_184 =>
            -- reg_a = a3_X; reg_b = a7_X; reg_acc = reg_o >> 272; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_185 =>
            -- reg_a = o3_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_186 =>
            -- reg_a = a4_X; reg_b = a6_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_187 =>
            -- reg_a = o4_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_188 =>
            -- reg_a = a5_X; reg_b = a5_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_189 =>
            -- reg_a = o5_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_190 =>
            -- reg_a = o6_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_191 =>
            -- reg_a = o7_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_192 =>
            -- reg_a = a4_X; reg_b = a7_X; reg_acc = reg_o >> 272; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_193 =>
            -- reg_a = o4_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_194 =>
            -- reg_a = a5_X; reg_b = a6_X; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_195 =>
            -- reg_a = o5_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_196 =>
            -- reg_a = o6_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_197 =>
            -- reg_a = o7_X; reg_b = primeSP4; reg_acc = reg_o; o3_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_198 =>
            -- reg_a = a5_X; reg_b = a7_X; reg_acc = reg_o >> 272; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_199 =>
            -- reg_a = o5_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_200 =>
            -- reg_a = a6_X; reg_b = a6_X; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_201 =>
            -- reg_a = o6_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_202 =>
            -- reg_a = o7_X; reg_b = primeSP5; reg_acc = reg_o; o4_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_203 =>
            -- reg_a = a6_X; reg_b = a7_X; reg_acc = reg_o >> 272; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_204 =>
            -- reg_a = o6_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_205 =>
            -- reg_a = o7_X; reg_b = primeSP6; reg_acc = reg_o; o5_X = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_206 =>
            -- reg_a = a7_X; reg_b = a7_X; reg_acc = reg_o >> 272; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_207 =>
            -- reg_a = o7_X; reg_b = primeSP7; reg_acc = reg_o; o6_X = reg_o; o7_X = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_direct_0 =>
            -- -- In case of size 1
            -- reg_a = a0_X; reg_b = b0_X; reg_acc = 0; o0_0 = reg_o; Enable sign a,b; operation : b +/- a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '1';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_direct_2 =>
            -- -- In case of size 2, 3, 4, 5, 6, 7, 8
            -- reg_a = a0_X; reg_b = b0_X; reg_acc = 0; o0_X = reg_o; operation : b +/- a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '1';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_direct_3 =>
            -- -- In case of size 2
            -- reg_a = a1_X; reg_b = b1_X; reg_acc = reg_o >> 272; o1_X = reg_o; Enable sign a, b; operation : b +/- a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '1';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_direct_5 =>
            -- -- In case of size 3, 4, 5, 6, 7, 8
            -- reg_a = a1_X; reg_b = b1_X; reg_acc = reg_o >> 272; o1_X = reg_o; operation : b +/- a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '1';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_direct_6 =>
            -- -- In case of size 3
            -- reg_a = a2_X; reg_b = b2_X; reg_acc = reg_o >> 272; o2_X = reg_o; Enable sign a,b; operation : b +/- a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '1';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_direct_8 =>
            -- -- In case of size 4, 5, 6, 7, 8
            -- reg_a = a2_X; reg_b = b2_X; reg_acc = reg_o >> 272; o2_X = reg_o; operation : b +/- a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '1';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_direct_9 =>
            -- -- In case of size 4
            -- reg_a = a3_X; reg_b = b3_X; reg_acc = reg_o >> 272; o3_X = reg_o; Enable sign a,b; operation : b +/- a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '1';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_direct_11 =>
            -- -- In case of size 4, 5, 6, 7, 8
            -- reg_a = a3_X; reg_b = b3_X; reg_acc = reg_o >> 272; o3_X = reg_o; operation : b +/- a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '1';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_direct_12 =>
            -- -- In case of size 5
            -- reg_a = a4_X; reg_b = b4_X; reg_acc = reg_o >> 272; o4_X = reg_o; Enable sign a,b; operation : b +/- a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '1';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_direct_14 =>
            -- -- In case of size 6, 7, 8
            -- reg_a = a4_X; reg_b = b4_X; reg_acc = reg_o >> 272; o4_X = reg_o; operation : b +/- a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '1';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_direct_15 =>
            -- -- In case of size 6
            -- reg_a = a5_X; reg_b = b5_X; reg_acc = reg_o >> 272; o5_X = reg_o; Enable sign a,b; operation : b +/- a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '1';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_direct_17 =>
            -- -- In case of size 7, 8
            -- reg_a = a5_X; reg_b = b5_X; reg_acc = reg_o >> 272; o5_X = reg_o; operation : b +/- a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '1';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_direct_18 =>
            -- -- In case of size 7
            -- reg_a = a6_X; reg_b = b6_X; reg_acc = reg_o >> 272; o6_X = reg_o; Enable sign a,b; operation : b +/- a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '1';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_direct_20 =>
            -- -- In case of size 8
            -- reg_a = a6_X; reg_b = b6_X; reg_acc = reg_o >> 272; o6_X = reg_o; operation : b +/- a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '1';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_direct_21 =>
            -- reg_a = a7_X; reg_b = b7_X; reg_acc = reg_o >> 272; o7_X = reg_o; Enable sign a,b; operation : b +/- a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "111";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '1';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_0 =>
            -- -- In case of size 1
            -- reg_a = a0_X; reg_b = 0; reg_acc = 0; Enable sign a,b; operation : b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '1';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_1 =>
            -- reg_a = 0; reg_b = prime0; reg_acc = reg_o; reg_s = reg_o_positive; Enable sign a,b; operation : -s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "11";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '1';
            next_mac_sel_reg_s_reg_o_sign <= '1';
            next_mac_reg_s_reg_o_positive <= '1';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_2 =>
            -- reg_a = 0; reg_b = prime0; reg_acc = reg_o; reg_s = reg_o_negative; Enable sign a,b; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "11";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '1';
            next_mac_sel_reg_s_reg_o_sign <= '1';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_3 =>
            -- reg_a = 0; reg_b = prime0; reg_acc = reg_o; o0_X = reg_o; reg_s = reg_o_negative; Enable sign a,b; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "11";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '1';
            next_mac_sel_reg_s_reg_o_sign <= '1';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_5 =>
            -- -- In case of size 2
            -- reg_a = a1_X; reg_b = 0; reg_acc = 0; Enable sign a,b; operation : b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '1';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_6 =>
            -- reg_a = a0_X; reg_b = prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_positive; operation : -s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '1';
            next_mac_sel_reg_s_reg_o_sign <= '1';
            next_mac_reg_s_reg_o_positive <= '1';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_7 =>
            -- reg_a = a1_X; reg_b = prime1; reg_acc = reg_o >> 272; o1_X = reg_o; Enable sign a,b; operation : -s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_8 =>
            -- reg_a = o0_X; reg_b = prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '1';
            next_mac_sel_reg_s_reg_o_sign <= '1';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_9 =>
            -- reg_a = o1_X; reg_b = prime1; reg_acc = reg_o >> 272; o1_X = reg_o; Enable sign a,b operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_10 =>
            -- reg_a = o0_X; reg_b = prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '1';
            next_mac_sel_reg_s_reg_o_sign <= '1';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_11 =>
            -- reg_a = o1_X; reg_b = prime1; reg_acc = reg_o >> 272; o1_X = reg_o; Enable sign a,b operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_13 =>
            -- -- In case of size 3
            -- reg_a = a2_X; reg_b = 0; reg_acc = 0; Enable sign a,b; operation : b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '1';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_14 =>
            -- reg_a = a0_X; reg_b = prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_positive; operation : -s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '1';
            next_mac_sel_reg_s_reg_o_sign <= '1';
            next_mac_reg_s_reg_o_positive <= '1';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_15 =>
            -- reg_a = a1_X; reg_b = prime1; reg_acc = reg_o >> 272; o1_X = reg_o; operation : -s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_16 =>
            -- reg_a = a2_X; reg_b = prime2; reg_acc = reg_o >> 272; o2_X = reg_o; Enable sign a,b; operation : -s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_17 =>
            -- reg_a = o0_X; reg_b = prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '1';
            next_mac_sel_reg_s_reg_o_sign <= '1';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_18 =>
            -- reg_a = o1_X; reg_b = prime1; reg_acc = reg_o >> 272; o1_X = reg_o; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_19 =>
            -- reg_a = o2_X; reg_b = prime2; reg_acc = reg_o >> 272; o2_X = reg_o; Enable sign a,b operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_20 =>
            -- reg_a = o0_X; reg_b = prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '1';
            next_mac_sel_reg_s_reg_o_sign <= '1';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_21 =>
            -- reg_a = o1_X; reg_b = prime1; reg_acc = reg_o >> 272; o1_X = reg_o; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_22 =>
            -- reg_a = o2_X; reg_b = prime2; reg_acc = reg_o >> 272; o2_X = reg_o; Enable sign a,b operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_24 =>
            -- -- In case of size 4
            -- reg_a = a3_X; reg_b = 0; reg_acc = 0; Enable sign a,b; operation : b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '1';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_25 =>
            -- reg_a = a0_X; reg_b = prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_positive; operation : -s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '1';
            next_mac_sel_reg_s_reg_o_sign <= '1';
            next_mac_reg_s_reg_o_positive <= '1';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_26 =>
            -- reg_a = a1_X; reg_b = prime1; reg_acc = reg_o >> 272; o1_X = reg_o; operation : -s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_27 =>
            -- reg_a = a2_X; reg_b = prime2; reg_acc = reg_o >> 272; o2_X = reg_o; operation : -s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_28 =>
            -- reg_a = a3_X; reg_b = prime3; reg_acc = reg_o >> 272; o3_X = reg_o; Enable sign a,b; operation : -s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_29 =>
            -- reg_a = o0_X; reg_b = prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '1';
            next_mac_sel_reg_s_reg_o_sign <= '1';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_30 =>
            -- reg_a = o1_X; reg_b = prime1; reg_acc = reg_o >> 272; o1_X = reg_o; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_31 =>
            -- reg_a = o2_X; reg_b = prime2; reg_acc = reg_o >> 272; o2_X = reg_o; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_32 =>
            -- reg_a = o3_X; reg_b = prime3; reg_acc = reg_o >> 272; o3_X = reg_o; Enable sign a,b; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_33 =>
            -- reg_a = o0_X; reg_b = prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '1';
            next_mac_sel_reg_s_reg_o_sign <= '1';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_34 =>
            -- reg_a = o1_X; reg_b = prime1; reg_acc = reg_o >> 272; o1_X = reg_o; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_35 =>
            -- reg_a = o2_X; reg_b = prime2; reg_acc = reg_o >> 272; o2_X = reg_o; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_36 =>
            -- reg_a = o3_X; reg_b = prime3; reg_acc = reg_o >> 272; o3_X = reg_o; Enable sign a,b; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_38 =>
            -- -- In case of size 5
            -- reg_a = a4_X; reg_b = 0; reg_acc = 0; Enable sign a,b; operation : b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '1';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_39 =>
            -- reg_a = a0_X; reg_b = prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_positive; operation : -s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '1';
            next_mac_sel_reg_s_reg_o_sign <= '1';
            next_mac_reg_s_reg_o_positive <= '1';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_40 =>
            -- reg_a = a1_X; reg_b = prime1; reg_acc = reg_o >> 272; o1_X = reg_o; operation : -s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_41 =>
            -- reg_a = a2_X; reg_b = prime2; reg_acc = reg_o >> 272; o2_X = reg_o; operation : -s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_42 =>
            -- reg_a = a3_X; reg_b = prime3; reg_acc = reg_o >> 272; o3_X = reg_o; operation : -s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_43 =>
            -- reg_a = a4_X; reg_b = prime4; reg_acc = reg_o >> 272; o4_X = reg_o; Enable sign a,b; operation : -s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_44 =>
            -- reg_a = o0_X; reg_b = prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '1';
            next_mac_sel_reg_s_reg_o_sign <= '1';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_45 =>
            -- reg_a = o1_X; reg_b = prime1; reg_acc = reg_o >> 272; o1_X = reg_o; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_46 =>
            -- reg_a = o2_X; reg_b = prime2; reg_acc = reg_o >> 272; o2_X = reg_o; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_47 =>
            -- reg_a = o3_X; reg_b = prime3; reg_acc = reg_o >> 272; o3_X = reg_o; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_48 =>
            -- reg_a = o4_X; reg_b = prime4; reg_acc = reg_o >> 272; o4_X = reg_o; Enable sign a,b; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_49 =>
            -- reg_a = o0_X; reg_b = prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '1';
            next_mac_sel_reg_s_reg_o_sign <= '1';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_50 =>
            -- reg_a = o1_X; reg_b = prime1; reg_acc = reg_o >> 272; o1_X = reg_o; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_51 =>
            -- reg_a = o2_X; reg_b = prime2; reg_acc = reg_o >> 272; o2_X = reg_o; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_52 =>
            -- reg_a = o3_X; reg_b = prime3; reg_acc = reg_o >> 272; o3_X = reg_o; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_53 =>
            -- reg_a = o4_X; reg_b = prime4; reg_acc = reg_o >> 272; o4_X = reg_o; Enable sign a,b; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_55 =>
            -- -- In case of size 6
            -- reg_a = a5_X; reg_b = 0; reg_acc = 0; Enable sign a,b; operation : b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '1';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_56 =>
            -- reg_a = a0_X; reg_b = prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_positive; operation : -s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '1';
            next_mac_sel_reg_s_reg_o_sign <= '1';
            next_mac_reg_s_reg_o_positive <= '1';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_57 =>
            -- reg_a = a1_X; reg_b = prime1; reg_acc = reg_o >> 272; o1_X = reg_o; operation : -s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_58 =>
            -- reg_a = a2_X; reg_b = prime2; reg_acc = reg_o >> 272; o2_X = reg_o; operation : -s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_59 =>
            -- reg_a = a3_X; reg_b = prime3; reg_acc = reg_o >> 272; o3_X = reg_o; operation : -s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_60 =>
            -- reg_a = a4_X; reg_b = prime4; reg_acc = reg_o >> 272; o4_X = reg_o; operation : -s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_61 =>
            -- reg_a = a5_X; reg_b = prime5; reg_acc = reg_o >> 272; o5_X = reg_o; Enable sign a,b; operation : -s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_62 =>
            -- reg_a = o0_X; reg_b = prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '1';
            next_mac_sel_reg_s_reg_o_sign <= '1';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_63 =>
            -- reg_a = o1_X; reg_b = prime1; reg_acc = reg_o >> 272; o1_X = reg_o; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_64 =>
            -- reg_a = o2_X; reg_b = prime2; reg_acc = reg_o >> 272; o2_X = reg_o; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_65 =>
            -- reg_a = o3_X; reg_b = prime3; reg_acc = reg_o >> 272; o3_X = reg_o; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_66 =>
            -- reg_a = o4_X; reg_b = prime4; reg_acc = reg_o >> 272; o4_X = reg_o; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_67 =>
            -- reg_a = o5_X; reg_b = prime5; reg_acc = reg_o >> 272; o5_X = reg_o; Enable sign a,b; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_68 =>
            -- reg_a = o0_X; reg_b = prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '1';
            next_mac_sel_reg_s_reg_o_sign <= '1';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_69 =>
            -- reg_a = o1_X; reg_b = prime1; reg_acc = reg_o >> 272; o1_X = reg_o; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_70 =>
            -- reg_a = o2_X; reg_b = prime2; reg_acc = reg_o >> 272; o2_X = reg_o; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_71 =>
            -- reg_a = o3_X; reg_b = prime3; reg_acc = reg_o >> 272; o3_X = reg_o; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_72 =>
            -- reg_a = o4_X; reg_b = prime4; reg_acc = reg_o >> 272; o4_X = reg_o; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_73 =>
            -- reg_a = o5_X; reg_b = prime5; reg_acc = reg_o >> 272; o5_X = reg_o; Enable sign a,b; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_75 =>
            -- -- In case of size 7
            -- reg_a = a6_X; reg_b = 0; reg_acc = 0; Enable sign a,b; operation : b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '1';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_76 =>
            -- reg_a = a0_X; reg_b = prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_positive; operation : -s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '1';
            next_mac_sel_reg_s_reg_o_sign <= '1';
            next_mac_reg_s_reg_o_positive <= '1';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_77 =>
            -- reg_a = a1_X; reg_b = prime1; reg_acc = reg_o >> 272; o1_X = reg_o; operation : -s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_78 =>
            -- reg_a = a2_X; reg_b = prime2; reg_acc = reg_o >> 272; o2_X = reg_o; operation : -s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_79 =>
            -- reg_a = a3_X; reg_b = prime3; reg_acc = reg_o >> 272; o3_X = reg_o; operation : -s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_80 =>
            -- reg_a = a4_X; reg_b = prime4; reg_acc = reg_o >> 272; o4_X = reg_o; operation : -s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_81 =>
            -- reg_a = a5_X; reg_b = prime5; reg_acc = reg_o >> 272; o5_X = reg_o; operation : -s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_82 =>
            -- reg_a = a6_X; reg_b = prime6; reg_acc = reg_o >> 272; o6_X = reg_o; Enable sign a,b; operation : -s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_83 =>
            -- reg_a = o0_X; reg_b = prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '1';
            next_mac_sel_reg_s_reg_o_sign <= '1';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_84 =>
            -- reg_a = o1_X; reg_b = prime1; reg_acc = reg_o >> 272; o1_X = reg_o; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_85 =>
            -- reg_a = o2_X; reg_b = prime2; reg_acc = reg_o >> 272; o2_X = reg_o; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_86 =>
            -- reg_a = o3_X; reg_b = prime3; reg_acc = reg_o >> 272; o3_X = reg_o; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_87 =>
            -- reg_a = o4_X; reg_b = prime4; reg_acc = reg_o >> 272; o4_X = reg_o; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_88 =>
            -- reg_a = o5_X; reg_b = prime5; reg_acc = reg_o >> 272; o5_X = reg_o; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_89 =>
            -- reg_a = o6_X; reg_b = prime6; reg_acc = reg_o >> 272; o6_X = reg_o; Enable sign a,b; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_90 =>
            -- reg_a = o0_X; reg_b = prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '1';
            next_mac_sel_reg_s_reg_o_sign <= '1';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_91 =>
            -- reg_a = o1_X; reg_b = prime1; reg_acc = reg_o >> 272; o1_X = reg_o; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_92 =>
            -- reg_a = o2_X; reg_b = prime2; reg_acc = reg_o >> 272; o2_X = reg_o; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_93 =>
            -- reg_a = o3_X; reg_b = prime3; reg_acc = reg_o >> 272; o3_X = reg_o; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_94 =>
            -- reg_a = o4_X; reg_b = prime4; reg_acc = reg_o >> 272; o4_X = reg_o; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_95 =>
            -- reg_a = o5_X; reg_b = prime5; reg_acc = reg_o >> 272; o5_X = reg_o; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_96 =>
            -- reg_a = o6_X; reg_b = prime6; reg_acc = reg_o >> 272; o6_X = reg_o; Enable sign a,b; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_98 =>
            -- -- In case of size 8
            -- reg_a = a7_X; reg_b = 0; reg_acc = 0; Enable sign a,b; operation : b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "111";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '1';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_99 =>
            -- reg_a = a0_X; reg_b = prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_positive; operation : -s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '1';
            next_mac_sel_reg_s_reg_o_sign <= '1';
            next_mac_reg_s_reg_o_positive <= '1';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_100 =>
            -- reg_a = a1_X; reg_b = prime1; reg_acc = reg_o >> 272; o1_X = reg_o; operation : -s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_101 =>
            -- reg_a = a2_X; reg_b = prime2; reg_acc = reg_o >> 272; o2_X = reg_o; operation : -s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_102 =>
            -- reg_a = a3_X; reg_b = prime3; reg_acc = reg_o >> 272; o3_X = reg_o; operation : -s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_103 =>
            -- reg_a = a4_X; reg_b = prime4; reg_acc = reg_o >> 272; o4_X = reg_o; operation : -s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_104 =>
            -- reg_a = a5_X; reg_b = prime5; reg_acc = reg_o >> 272; o5_X = reg_o; operation : -s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_105 =>
            -- reg_a = a6_X; reg_b = prime6; reg_acc = reg_o >> 272; o6_X = reg_o; operation : -s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_106 =>
            -- reg_a = a7_X; reg_b = prime7; reg_acc = reg_o >> 272; o7_X = reg_o; Enable sign a,b; operation : -s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "111";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_107 =>
            -- reg_a = o0_X; reg_b = prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '1';
            next_mac_sel_reg_s_reg_o_sign <= '1';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_108 =>
            -- reg_a = o1_X; reg_b = prime1; reg_acc = reg_o >> 272; o1_X = reg_o; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_109 =>
            -- reg_a = o2_X; reg_b = prime2; reg_acc = reg_o >> 272; o2_X = reg_o; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_110 =>
            -- reg_a = o3_X; reg_b = prime3; reg_acc = reg_o >> 272; o3_X = reg_o; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_111 =>
            -- reg_a = o4_X; reg_b = prime4; reg_acc = reg_o >> 272; o4_X = reg_o; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_112 =>
            -- reg_a = o5_X; reg_b = prime5; reg_acc = reg_o >> 272; o5_X = reg_o; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_113 =>
            -- reg_a = o6_X; reg_b = prime6; reg_acc = reg_o >> 272; o6_X = reg_o; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_114 =>
            -- reg_a = o7_X; reg_b = prime7; reg_acc = reg_o >> 272; o7_X = reg_o; Enable sign a,b; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "111";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_115 =>
            -- reg_a = o0_X; reg_b = prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '1';
            next_mac_sel_reg_s_reg_o_sign <= '1';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_116 =>
            -- reg_a = o1_X; reg_b = prime1; reg_acc = reg_o >> 272; o1_X = reg_o; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "001";
            next_sm_specific_mac_address_b <= "001";
            next_sm_specific_mac_address_o <= "001";
            next_sm_specific_mac_next_address_o <= "010";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_117 =>
            -- reg_a = o2_X; reg_b = prime2; reg_acc = reg_o >> 272; o2_X = reg_o; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "010";
            next_sm_specific_mac_address_b <= "010";
            next_sm_specific_mac_address_o <= "010";
            next_sm_specific_mac_next_address_o <= "011";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_118 =>
            -- reg_a = o3_X; reg_b = prime3; reg_acc = reg_o >> 272; o3_X = reg_o; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "011";
            next_sm_specific_mac_address_b <= "011";
            next_sm_specific_mac_address_o <= "011";
            next_sm_specific_mac_next_address_o <= "100";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_119 =>
            -- reg_a = o4_X; reg_b = prime4; reg_acc = reg_o >> 272; o4_X = reg_o; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "100";
            next_sm_specific_mac_address_b <= "100";
            next_sm_specific_mac_address_o <= "100";
            next_sm_specific_mac_next_address_o <= "101";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_120 =>
            -- reg_a = o5_X; reg_b = prime5; reg_acc = reg_o >> 272; o5_X = reg_o; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "101";
            next_sm_specific_mac_address_b <= "101";
            next_sm_specific_mac_address_o <= "101";
            next_sm_specific_mac_next_address_o <= "110";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_121 =>
            -- reg_a = o6_X; reg_b = prime6; reg_acc = reg_o >> 272; o6_X = reg_o; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "110";
            next_sm_specific_mac_address_b <= "110";
            next_sm_specific_mac_address_o <= "110";
            next_sm_specific_mac_next_address_o <= "111";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_122 =>
            -- reg_a = o7_X; reg_b = prime7; reg_acc = reg_o >> 272; o7_X = reg_o; Enable sign a,b; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "111";
            next_sm_specific_mac_address_b <= "111";
            next_sm_specific_mac_address_o <= "111";
            next_sm_specific_mac_next_address_o <= "000";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when nop_4_stages =>
        -- reg_a = 0; reg_b = 0; reg_acc = 0; operation : b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "11";
            next_mac_clear_reg_b <= '1';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when nop_8_stages =>
        -- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "000";
            next_sm_specific_mac_address_b <= "000";
            next_sm_specific_mac_address_o <= "000";
            next_sm_specific_mac_next_address_o <= "001";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "11";
            next_mac_clear_reg_b <= '1';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
--        when others => 
--            next_sm_free_flag <= '0';
--            next_sm_rotation_size <= "11";
--            next_sm_circular_shift_enable <= '0';
--            next_sel_address_a <= '0';
--            next_sel_address_b_prime <= "00";
--            next_sm_specific_mac_address_a <= "000";
--            next_sm_specific_mac_address_b <= "000";
--            next_sm_specific_mac_address_o <= "000";
--            next_sm_specific_mac_next_address_o <= "001";
--            next_mac_enable_signed_a <= '0';
--            next_mac_enable_signed_b <= '0';
--            next_mac_sel_load_reg_a <= "11";
--            next_mac_clear_reg_b <= '1';
--            next_mac_clear_reg_acc <= '1';
--            next_mac_sel_shift_reg_o <= '0';
--            next_mac_enable_update_reg_s <= '0';
--            next_mac_sel_reg_s_reg_o_sign <= '0';
--            next_mac_reg_s_reg_o_positive <= '0';
--            next_sm_sign_a_mode <= '0';
--            next_sm_mac_operation_mode <= "10";
--            next_mac_enable_reg_s_mask <= '0';
--            next_mac_subtraction_reg_a_b <= '0';
--            next_mac_sel_multiply_two_a_b <= '0';
--            next_mac_sel_reg_y_output <= '0';
--            next_sm_mac_write_enable_output <= '0';
--            next_mac_memory_double_mode <= '0';
--            next_mac_memory_only_write_mode <= '0';
--            next_base_address_generator_o_increment_previous_address <= '0';
    end case;
end process;

update_state : process(actual_state, instruction_values_valid, instruction_type, prime_line_equal_one, operands_size, penultimate_operation)
begin
case (actual_state) is
        when reset =>
            next_state <= decode_instruction;
        when decode_instruction =>
            next_state <= decode_instruction;
            if(instruction_values_valid = '1') then
                if(instruction_type = "0000") then
                    if(operands_size = "000") then
                        next_state <= multiplication_direct_0;
                    else
                        next_state <= multiplication_direct_2;
                    end if;
                elsif(instruction_type = "0001") then
                    if(operands_size = "000") then
                        next_state <= square_direct_0;
                    else
                        next_state <= square_direct_2;
                    end if;
                elsif(instruction_type = "0010") then
                    if(prime_line_equal_one = '1') then
                        case (operands_size) is
                            when "000" =>
                                next_state <= multiplication_with_reduction_special_prime_0;
                            when "001"| "010"| "011" =>
                                next_state <= multiplication_with_reduction_special_prime_3;
                            when "100"| "101" =>
                                next_state <= multiplication_with_reduction_special_prime_47;
                            when others => 
                                next_state <= multiplication_with_reduction_special_prime_130;
                        end case;
                    else
                        if(operands_size = "000") then
                            next_state <= multiplication_with_reduction_0;
                        else
                            next_state <= multiplication_with_reduction_5;
                        end if;
                    end if;
                elsif(instruction_type = "0011") then
                    if(prime_line_equal_one = '1') then
                        case (operands_size) is
                            when "000" =>
                                next_state <= square_with_reduction_special_prime_0;
                            when "001"| "010"| "011" =>
                                next_state <= square_with_reduction_special_prime_3;
                            when "100"| "101" =>
                                next_state <= square_with_reduction_special_prime_37;
                            when others => 
                                next_state <= square_with_reduction_special_prime_100;
                        end case;
                    else
                        if(operands_size = "000") then
                            next_state <= square_with_reduction_0;
                        else
                            next_state <= square_with_reduction_5;
                        end if;
                    end if;
                elsif(instruction_type = "0100") then
                    if(operands_size = "000") then
                        next_state <= addition_subtraction_direct_0;
                    else
                        next_state <= addition_subtraction_direct_2;
                    end if;
                elsif(instruction_type = "0101") then
                    if(operands_size = "000") then
                        next_state <= iterative_modular_reduction_0;
                    elsif(operands_size = "001") then
                        next_state <= iterative_modular_reduction_5;
                    elsif(operands_size = "010") then
                        next_state <= iterative_modular_reduction_13;
                    elsif(operands_size = "011") then
                        next_state <= iterative_modular_reduction_24;
                    elsif(operands_size = "100") then
                        next_state <= iterative_modular_reduction_38;
                    elsif(operands_size = "101") then
                        next_state <= iterative_modular_reduction_55;
                    elsif(operands_size = "110") then
                        next_state <= iterative_modular_reduction_75;
                    else
                        next_state <= iterative_modular_reduction_98;
                    end if;
                end if;
            end if;
        when multiplication_direct_0 =>
            next_state <= multiplication_direct_0;
            if(penultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when multiplication_direct_2 =>
            next_state <= multiplication_direct_2;
            if(penultimate_operation = '1') then
                if(operands_size = "001") then
                    next_state <= multiplication_direct_3;
                else
                    next_state <= multiplication_direct_7;
                end if;
            end if;
        when multiplication_direct_3 =>
            next_state <= multiplication_direct_3;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_4;
            end if;
        when multiplication_direct_4 =>
            next_state <= multiplication_direct_4;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_5;
            end if;
        when multiplication_direct_5 =>
            next_state <= multiplication_direct_5;
            if(penultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when multiplication_direct_7 =>
            next_state <= multiplication_direct_7;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_8;
            end if;
        when multiplication_direct_8 =>
            next_state <= multiplication_direct_8;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_9;
            end if;
        when multiplication_direct_9 =>
            next_state <= multiplication_direct_9;
            if(penultimate_operation = '1') then
                if(operands_size = "010") then
                    next_state <= multiplication_direct_10;
                else
                    next_state <= multiplication_direct_16;
                end if;
            end if;
        when multiplication_direct_10 =>
            next_state <= multiplication_direct_10;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_11;
            end if;
        when multiplication_direct_11 =>
            next_state <= multiplication_direct_11;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_12;
            end if;
        when multiplication_direct_12 =>
            next_state <= multiplication_direct_12;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_13;
            end if;
        when multiplication_direct_13 =>
            next_state <= multiplication_direct_13;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_14;
            end if;
        when multiplication_direct_14 =>
            next_state <= multiplication_direct_14;
            if(penultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when multiplication_direct_16 =>
            next_state <= multiplication_direct_16;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_17;
            end if;
        when multiplication_direct_17 =>
            next_state <= multiplication_direct_17;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_18;
            end if;
        when multiplication_direct_18 =>
            next_state <= multiplication_direct_18;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_19;
            end if;
        when multiplication_direct_19 =>
            next_state <= multiplication_direct_19;
            if(penultimate_operation = '1') then
                if(operands_size = "011") then
                    next_state <= multiplication_direct_20;
                else
                    next_state <= multiplication_direct_29;
                end if;
            end if;
        when multiplication_direct_20 =>
            next_state <= multiplication_direct_20;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_21;
            end if;
        when multiplication_direct_21 =>
            next_state <= multiplication_direct_21;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_22;
            end if;
        when multiplication_direct_22 =>
            next_state <= multiplication_direct_22;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_23;
            end if;
        when multiplication_direct_23 =>
            next_state <= multiplication_direct_23;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_24;
            end if;
        when multiplication_direct_24 =>
            next_state <= multiplication_direct_24;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_25;
            end if;
        when multiplication_direct_25 =>
            next_state <= multiplication_direct_25;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_26;
            end if;
        when multiplication_direct_26 =>
            next_state <= multiplication_direct_26;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_27;
            end if;
        when multiplication_direct_27 =>
            next_state <= multiplication_direct_27;
            if(penultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when multiplication_direct_29 =>
            next_state <= multiplication_direct_29;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_30;
            end if;
        when multiplication_direct_30 =>
            next_state <= multiplication_direct_30;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_31;
            end if;
        when multiplication_direct_31 =>
            next_state <= multiplication_direct_31;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_32;
            end if;
        when multiplication_direct_32 =>
            next_state <= multiplication_direct_32;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_33;
            end if;
        when multiplication_direct_33 =>
            next_state <= multiplication_direct_33;
            if(penultimate_operation = '1') then
                if(operands_size = "100") then
                    next_state <= multiplication_direct_34;
                else
                    next_state <= multiplication_direct_47;
                end if;
            end if;
        when multiplication_direct_34 =>
            next_state <= multiplication_direct_34;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_35;
            end if;
        when multiplication_direct_35 =>
            next_state <= multiplication_direct_35;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_36;
            end if;
        when multiplication_direct_36 =>
            next_state <= multiplication_direct_36;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_37;
            end if;
        when multiplication_direct_37 =>
            next_state <= multiplication_direct_37;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_38;
            end if;
        when multiplication_direct_38 =>
            next_state <= multiplication_direct_38;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_39;
            end if;
        when multiplication_direct_39 =>
            next_state <= multiplication_direct_39;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_40;
            end if;
        when multiplication_direct_40 =>
            next_state <= multiplication_direct_40;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_41;
            end if;
        when multiplication_direct_41 =>
            next_state <= multiplication_direct_41;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_42;
            end if;
        when multiplication_direct_42 =>
            next_state <= multiplication_direct_42;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_43;
            end if;
        when multiplication_direct_43 =>
            next_state <= multiplication_direct_43;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_44;
            end if;
        when multiplication_direct_44 =>
            next_state <= multiplication_direct_44;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_45;
            end if;
        when multiplication_direct_45 =>
            next_state <= multiplication_direct_45;
            if(penultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when multiplication_direct_47 =>
            next_state <= multiplication_direct_47;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_48;
            end if;
        when multiplication_direct_48 =>
            next_state <= multiplication_direct_48;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_49;
            end if;
        when multiplication_direct_49 =>
            next_state <= multiplication_direct_49;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_50;
            end if;
        when multiplication_direct_50 =>
            next_state <= multiplication_direct_50;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_51;
            end if;
        when multiplication_direct_51 =>
            next_state <= multiplication_direct_51;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_52;
            end if;
        when multiplication_direct_52 =>
            next_state <= multiplication_direct_52;
            if(penultimate_operation = '1') then
                if(operands_size = "101") then
                    next_state <= multiplication_direct_53;
                else
                    next_state <= multiplication_direct_71;
                end if;
            end if;
        when multiplication_direct_53 =>
            next_state <= multiplication_direct_53;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_54;
            end if;
        when multiplication_direct_54 =>
            next_state <= multiplication_direct_54;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_55;
            end if;
        when multiplication_direct_55 =>
            next_state <= multiplication_direct_55;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_56;
            end if;
        when multiplication_direct_56 =>
            next_state <= multiplication_direct_56;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_57;
            end if;
        when multiplication_direct_57 =>
            next_state <= multiplication_direct_57;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_58;
            end if;
        when multiplication_direct_58 =>
            next_state <= multiplication_direct_58;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_59;
            end if;
        when multiplication_direct_59 =>
            next_state <= multiplication_direct_59;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_60;
            end if;
        when multiplication_direct_60 =>
            next_state <= multiplication_direct_60;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_61;
            end if;
        when multiplication_direct_61 =>
            next_state <= multiplication_direct_61;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_62;
            end if;
        when multiplication_direct_62 =>
            next_state <= multiplication_direct_62;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_63;
            end if;
        when multiplication_direct_63 =>
            next_state <= multiplication_direct_63;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_64;
            end if;
        when multiplication_direct_64 =>
            next_state <= multiplication_direct_64;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_65;
            end if;
        when multiplication_direct_65 =>
            next_state <= multiplication_direct_65;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_66;
            end if;
        when multiplication_direct_66 =>
            next_state <= multiplication_direct_66;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_67;
            end if;
        when multiplication_direct_67 =>
            next_state <= multiplication_direct_67;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_68;
            end if;
        when multiplication_direct_68 =>
            next_state <= multiplication_direct_68;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_69;
            end if;
        when multiplication_direct_69 =>
            next_state <= multiplication_direct_69;
            if(penultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when multiplication_direct_71 =>
            next_state <= multiplication_direct_71;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_72;
            end if;
        when multiplication_direct_72 =>
            next_state <= multiplication_direct_72;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_73;
            end if;
        when multiplication_direct_73 =>
            next_state <= multiplication_direct_73;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_74;
            end if;
        when multiplication_direct_74 =>
            next_state <= multiplication_direct_74;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_75;
            end if;
        when multiplication_direct_75 =>
            next_state <= multiplication_direct_75;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_76;
            end if;
        when multiplication_direct_76 =>
            next_state <= multiplication_direct_76;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_77;
            end if;
        when multiplication_direct_77 =>
            next_state <= multiplication_direct_77;
            if(penultimate_operation = '1') then
                if(operands_size = "110") then
                    next_state <= multiplication_direct_78;
                else
                    next_state <= multiplication_direct_102;
                end if;
            end if;
        when multiplication_direct_78 =>
            next_state <= multiplication_direct_78;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_79;
            end if;
        when multiplication_direct_79 =>
            next_state <= multiplication_direct_79;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_80;
            end if;
        when multiplication_direct_80 =>
            next_state <= multiplication_direct_80;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_81;
            end if;
        when multiplication_direct_81 =>
            next_state <= multiplication_direct_81;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_82;
            end if;
        when multiplication_direct_82 =>
            next_state <= multiplication_direct_82;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_83;
            end if;
        when multiplication_direct_83 =>
            next_state <= multiplication_direct_83;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_84;
            end if;
        when multiplication_direct_84 =>
            next_state <= multiplication_direct_84;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_85;
            end if;
        when multiplication_direct_85 =>
            next_state <= multiplication_direct_85;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_86;
            end if;
        when multiplication_direct_86 =>
            next_state <= multiplication_direct_86;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_87;
            end if;
        when multiplication_direct_87 =>
            next_state <= multiplication_direct_87;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_88;
            end if;
        when multiplication_direct_88 =>
            next_state <= multiplication_direct_88;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_89;
            end if;
        when multiplication_direct_89 =>
            next_state <= multiplication_direct_89;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_90;
            end if;
        when multiplication_direct_90 =>
            next_state <= multiplication_direct_90;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_91;
            end if;
        when multiplication_direct_91 =>
            next_state <= multiplication_direct_91;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_92;
            end if;
        when multiplication_direct_92 =>
            next_state <= multiplication_direct_92;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_93;
            end if;
        when multiplication_direct_93 =>
            next_state <= multiplication_direct_93;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_94;
            end if;
        when multiplication_direct_94 =>
            next_state <= multiplication_direct_94;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_95;
            end if;
        when multiplication_direct_95 =>
            next_state <= multiplication_direct_95;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_96;
            end if;
        when multiplication_direct_96 =>
            next_state <= multiplication_direct_96;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_97;
            end if;
        when multiplication_direct_97 =>
            next_state <= multiplication_direct_97;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_98;
            end if;
        when multiplication_direct_98 =>
            next_state <= multiplication_direct_98;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_99;
            end if;
        when multiplication_direct_99 =>
            next_state <= multiplication_direct_99;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_100;
            end if;
        when multiplication_direct_100 =>
            next_state <= multiplication_direct_100;
            if(penultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when multiplication_direct_102 =>
            next_state <= multiplication_direct_102;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_103;
            end if;
        when multiplication_direct_103 =>
            next_state <= multiplication_direct_103;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_104;
            end if;
        when multiplication_direct_104 =>
            next_state <= multiplication_direct_104;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_105;
            end if;
        when multiplication_direct_105 =>
            next_state <= multiplication_direct_105;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_106;
            end if;
        when multiplication_direct_106 =>
            next_state <= multiplication_direct_106;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_107;
            end if;
        when multiplication_direct_107 =>
            next_state <= multiplication_direct_107;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_108;
            end if;
        when multiplication_direct_108 =>
            next_state <= multiplication_direct_108;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_109;
            end if;
        when multiplication_direct_109 =>
            next_state <= multiplication_direct_109;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_110;
            end if;
        when multiplication_direct_110 =>
            next_state <= multiplication_direct_110;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_111;
            end if;
        when multiplication_direct_111 =>
            next_state <= multiplication_direct_111;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_112;
            end if;
        when multiplication_direct_112 =>
            next_state <= multiplication_direct_112;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_113;
            end if;
        when multiplication_direct_113 =>
            next_state <= multiplication_direct_113;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_114;
            end if;
        when multiplication_direct_114 =>
            next_state <= multiplication_direct_114;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_115;
            end if;
        when multiplication_direct_115 =>
            next_state <= multiplication_direct_115;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_116;
            end if;
        when multiplication_direct_116 =>
            next_state <= multiplication_direct_116;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_117;
            end if;
        when multiplication_direct_117 =>
            next_state <= multiplication_direct_117;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_118;
            end if;
        when multiplication_direct_118 =>
            next_state <= multiplication_direct_118;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_119;
            end if;
        when multiplication_direct_119 =>
            next_state <= multiplication_direct_119;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_120;
            end if;
        when multiplication_direct_120 =>
            next_state <= multiplication_direct_120;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_121;
            end if;
        when multiplication_direct_121 =>
            next_state <= multiplication_direct_121;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_122;
            end if;
        when multiplication_direct_122 =>
            next_state <= multiplication_direct_122;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_123;
            end if;
        when multiplication_direct_123 =>
            next_state <= multiplication_direct_123;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_124;
            end if;
        when multiplication_direct_124 =>
            next_state <= multiplication_direct_124;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_125;
            end if;
        when multiplication_direct_125 =>
            next_state <= multiplication_direct_125;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_126;
            end if;
        when multiplication_direct_126 =>
            next_state <= multiplication_direct_126;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_127;
            end if;
        when multiplication_direct_127 =>
            next_state <= multiplication_direct_127;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_128;
            end if;
        when multiplication_direct_128 =>
            next_state <= multiplication_direct_128;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_129;
            end if;
        when multiplication_direct_129 =>
            next_state <= multiplication_direct_129;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_130;
            end if;
        when multiplication_direct_130 =>
            next_state <= multiplication_direct_130;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_131;
            end if;
        when multiplication_direct_131 =>
            next_state <= multiplication_direct_131;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_132;
            end if;
        when multiplication_direct_132 =>
            next_state <= multiplication_direct_132;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_133;
            end if;
        when multiplication_direct_133 =>
            next_state <= multiplication_direct_133;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_134;
            end if;
        when multiplication_direct_134 =>
            next_state <= multiplication_direct_134;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_135;
            end if;
        when multiplication_direct_135 =>
            next_state <= multiplication_direct_135;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_136;
            end if;
        when multiplication_direct_136 =>
            next_state <= multiplication_direct_136;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_137;
            end if;
        when multiplication_direct_137 =>
            next_state <= multiplication_direct_137;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_138;
            end if;
        when multiplication_direct_138 =>
            next_state <= multiplication_direct_138;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_139;
            end if;
        when multiplication_direct_139 =>
            next_state <= multiplication_direct_139;
            if(penultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when square_direct_0 => 
            next_state <= square_direct_0;
            if(penultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when square_direct_2 => 
            next_state <= square_direct_2;
            if(penultimate_operation = '1') then
                if(operands_size = "001") then
                    next_state <= square_direct_3;
                else
                    next_state <= square_direct_6;
                end if;
            end if;
        when square_direct_3 => 
            next_state <= square_direct_3;
            if(penultimate_operation = '1') then
                next_state <= square_direct_4;
            end if;
        when square_direct_4 => 
            next_state <= square_direct_4;
            if(penultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when square_direct_6 => 
            next_state <= square_direct_6;
            if(penultimate_operation = '1') then
                next_state <= square_direct_7;
            end if;
        when square_direct_7 => 
            next_state <= square_direct_7;
            if(penultimate_operation = '1') then
                if(operands_size = "010") then
                    next_state <= square_direct_8;
                else
                    next_state <= square_direct_12;
                end if;
            end if;
        when square_direct_8 => 
            next_state <= square_direct_8;
            if(penultimate_operation = '1') then
                next_state <= square_direct_9;
            end if;
        when square_direct_9 => 
            next_state <= square_direct_9;
            if(penultimate_operation = '1') then
                next_state <= square_direct_10;
            end if;
        when square_direct_10 => 
            next_state <= square_direct_10;
            if(penultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when square_direct_12 => 
            next_state <= square_direct_12;
            if(penultimate_operation = '1') then
                next_state <= square_direct_13;
            end if;
        when square_direct_13 => 
            next_state <= square_direct_13;
            if(penultimate_operation = '1') then
                if(operands_size = "011") then
                    next_state <= square_direct_14;
                else
                    next_state <= square_direct_20;
                end if;
            end if;
        when square_direct_14 => 
            next_state <= square_direct_14;
            if(penultimate_operation = '1') then
                next_state <= square_direct_15;
            end if;
        when square_direct_15 => 
            next_state <= square_direct_15;
            if(penultimate_operation = '1') then
                next_state <= square_direct_16;
            end if;
        when square_direct_16 => 
            next_state <= square_direct_16;
            if(penultimate_operation = '1') then
                next_state <= square_direct_17;
            end if;
        when square_direct_17 => 
            next_state <= square_direct_17;
            if(penultimate_operation = '1') then
                next_state <= square_direct_18;
            end if;
        when square_direct_18 => 
            next_state <= square_direct_18;
            if(penultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when square_direct_20 => 
            next_state <= square_direct_20;
            if(penultimate_operation = '1') then
                next_state <= square_direct_21;
            end if;
        when square_direct_21 => 
            next_state <= square_direct_21;
            if(penultimate_operation = '1') then
                next_state <= square_direct_22;
            end if;
        when square_direct_22 => 
            next_state <= square_direct_22;
            if(penultimate_operation = '1') then
                if(operands_size = "100") then
                    next_state <= square_direct_23;
                else
                    next_state <= square_direct_31;
                end if;
            end if;
        when square_direct_23 => 
            next_state <= square_direct_23;
            if(penultimate_operation = '1') then
                next_state <= square_direct_24;
            end if;
        when square_direct_24 => 
            next_state <= square_direct_24;
            if(penultimate_operation = '1') then
                next_state <= square_direct_25;
            end if;
        when square_direct_25 => 
            next_state <= square_direct_25;
            if(penultimate_operation = '1') then
                next_state <= square_direct_26;
            end if;
        when square_direct_26 => 
            next_state <= square_direct_26;
            if(penultimate_operation = '1') then
                next_state <= square_direct_27;
            end if;
        when square_direct_27 => 
            next_state <= square_direct_27;
            if(penultimate_operation = '1') then
                next_state <= square_direct_28;
            end if;
        when square_direct_28 => 
            next_state <= square_direct_28;
            if(penultimate_operation = '1') then
                next_state <= square_direct_29;
            end if;
        when square_direct_29 => 
            next_state <= square_direct_29;
            if(penultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when square_direct_31 => 
            next_state <= square_direct_31;
            if(penultimate_operation = '1') then
                next_state <= square_direct_32;
            end if;
        when square_direct_32 => 
            next_state <= square_direct_32;
            if(penultimate_operation = '1') then
                next_state <= square_direct_33;
            end if;
        when square_direct_33 => 
            next_state <= square_direct_33;
            if(penultimate_operation = '1') then
                if(operands_size = "101") then
                    next_state <= square_direct_34;
                else
                    next_state <= square_direct_45;
                end if;
            end if;
        when square_direct_34 => 
            next_state <= square_direct_34;
            if(penultimate_operation = '1') then
                next_state <= square_direct_35;
            end if;
        when square_direct_35 => 
            next_state <= square_direct_35;
            if(penultimate_operation = '1') then
                next_state <= square_direct_36;
            end if;
        when square_direct_36 => 
            next_state <= square_direct_36;
            if(penultimate_operation = '1') then
                next_state <= square_direct_37;
            end if;
        when square_direct_37 => 
            next_state <= square_direct_37;
            if(penultimate_operation = '1') then
                next_state <= square_direct_38;
            end if;
        when square_direct_38 => 
            next_state <= square_direct_38;
            if(penultimate_operation = '1') then
                next_state <= square_direct_39;
            end if;
        when square_direct_39 => 
            next_state <= square_direct_39;
            if(penultimate_operation = '1') then
                next_state <= square_direct_40;
            end if;
        when square_direct_40 => 
            next_state <= square_direct_40;
            if(penultimate_operation = '1') then
                next_state <= square_direct_41;
            end if;
        when square_direct_41 => 
            next_state <= square_direct_41;
            if(penultimate_operation = '1') then
                next_state <= square_direct_42;
            end if;
        when square_direct_42 => 
            next_state <= square_direct_42;
            if(penultimate_operation = '1') then
                next_state <= square_direct_43;
            end if;
        when square_direct_43 => 
            next_state <= square_direct_43;
            if(penultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when square_direct_45 => 
            next_state <= square_direct_45;
            if(penultimate_operation = '1') then
                next_state <= square_direct_46;
            end if;
        when square_direct_46 => 
            next_state <= square_direct_46;
            if(penultimate_operation = '1') then
                next_state <= square_direct_47;
            end if;
        when square_direct_47 => 
            next_state <= square_direct_47;
            if(penultimate_operation = '1') then
                next_state <= square_direct_48;
            end if;
        when square_direct_48 => 
            next_state <= square_direct_48;
            if(penultimate_operation = '1') then
                if(operands_size = "110") then
                    next_state <= square_direct_49;
                else
                    next_state <= square_direct_63;
                end if;
            end if;
        when square_direct_49 => 
            next_state <= square_direct_49;
            if(penultimate_operation = '1') then
                next_state <= square_direct_50;
            end if;
        when square_direct_50 => 
            next_state <= square_direct_50;
            if(penultimate_operation = '1') then
                next_state <= square_direct_51;
            end if;
        when square_direct_51 => 
            next_state <= square_direct_51;
            if(penultimate_operation = '1') then
                next_state <= square_direct_52;
            end if;
        when square_direct_52 => 
            next_state <= square_direct_52;
            if(penultimate_operation = '1') then
                next_state <= square_direct_53;
            end if;
        when square_direct_53 => 
            next_state <= square_direct_53;
            if(penultimate_operation = '1') then
                next_state <= square_direct_54;
            end if;
        when square_direct_54 => 
            next_state <= square_direct_54;
            if(penultimate_operation = '1') then
                next_state <= square_direct_55;
            end if;
        when square_direct_55 => 
            next_state <= square_direct_55;
            if(penultimate_operation = '1') then
                next_state <= square_direct_56;
            end if;
        when square_direct_56 => 
            next_state <= square_direct_56;
            if(penultimate_operation = '1') then
                next_state <= square_direct_57;
            end if;
        when square_direct_57 => 
            next_state <= square_direct_57;
            if(penultimate_operation = '1') then
                next_state <= square_direct_58;
            end if;
        when square_direct_58 => 
            next_state <= square_direct_58;
            if(penultimate_operation = '1') then
                next_state <= square_direct_59;
            end if;
        when square_direct_59 => 
            next_state <= square_direct_59;
            if(penultimate_operation = '1') then
                next_state <= square_direct_60;
            end if;
        when square_direct_60 => 
            next_state <= square_direct_60;
            if(penultimate_operation = '1') then
                next_state <= square_direct_61;
            end if;
        when square_direct_61 => 
            next_state <= square_direct_61;
            if(penultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when square_direct_63 => 
            next_state <= square_direct_63;
            if(penultimate_operation = '1') then
                next_state <= square_direct_64;
            end if;
        when square_direct_64 => 
            next_state <= square_direct_64;
            if(penultimate_operation = '1') then
                next_state <= square_direct_65;
            end if;
        when square_direct_65 => 
            next_state <= square_direct_65;
            if(penultimate_operation = '1') then
                next_state <= square_direct_66;
            end if;
        when square_direct_66 => 
            next_state <= square_direct_66;
            if(penultimate_operation = '1') then
                next_state <= square_direct_67;
            end if;
        when square_direct_67 => 
            next_state <= square_direct_67;
            if(penultimate_operation = '1') then
                next_state <= square_direct_68;
            end if;
        when square_direct_68 => 
            next_state <= square_direct_68;
            if(penultimate_operation = '1') then
                next_state <= square_direct_69;
            end if;
        when square_direct_69 => 
            next_state <= square_direct_69;
            if(penultimate_operation = '1') then
                next_state <= square_direct_70;
            end if;
        when square_direct_70 => 
            next_state <= square_direct_70;
            if(penultimate_operation = '1') then
                next_state <= square_direct_71;
            end if;
        when square_direct_71 => 
            next_state <= square_direct_71;
            if(penultimate_operation = '1') then
                next_state <= square_direct_72;
            end if;
        when square_direct_72 => 
            next_state <= square_direct_72;
            if(penultimate_operation = '1') then
                next_state <= square_direct_73;
            end if;
        when square_direct_73 => 
            next_state <= square_direct_73;
            if(penultimate_operation = '1') then
                next_state <= square_direct_74;
            end if;
        when square_direct_74 => 
            next_state <= square_direct_74;
            if(penultimate_operation = '1') then
                next_state <= square_direct_75;
            end if;
        when square_direct_75 => 
            next_state <= square_direct_75;
            if(penultimate_operation = '1') then
                next_state <= square_direct_76;
            end if;
        when square_direct_76 => 
            next_state <= square_direct_76;
            if(penultimate_operation = '1') then
                next_state <= square_direct_77;
            end if;
        when square_direct_77 => 
            next_state <= square_direct_77;
            if(penultimate_operation = '1') then
                next_state <= square_direct_78;
            end if;
        when square_direct_78 => 
            next_state <= square_direct_78;
            if(penultimate_operation = '1') then
                next_state <= square_direct_79;
            end if;
        when square_direct_79 => 
            next_state <= square_direct_79;
            if(penultimate_operation = '1') then
                next_state <= square_direct_80;
            end if;
        when square_direct_80 => 
            next_state <= square_direct_80;
            if(penultimate_operation = '1') then
                next_state <= square_direct_81;
            end if;
        when square_direct_81 => 
            next_state <= square_direct_81;
            if(penultimate_operation = '1') then
                next_state <= square_direct_82;
            end if;
        when square_direct_82 => 
            next_state <= square_direct_82;
            if(penultimate_operation = '1') then
                next_state <= square_direct_83;
            end if;
        when square_direct_83 => 
            next_state <= square_direct_83;
            if(penultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when multiplication_with_reduction_0 => 
            next_state <= multiplication_with_reduction_0;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_1;
            end if;
        when multiplication_with_reduction_1 => 
            next_state <= multiplication_with_reduction_1;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_2;
            end if;
        when multiplication_with_reduction_2 => 
            next_state <= multiplication_with_reduction_2;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_3;
            end if;
        when multiplication_with_reduction_3 => 
            next_state <= multiplication_with_reduction_3;
            if(penultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when multiplication_with_reduction_5 => 
            next_state <= multiplication_with_reduction_5;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_6;
            end if;
        when multiplication_with_reduction_6 => 
            next_state <= multiplication_with_reduction_6;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_7;
            end if;
        when multiplication_with_reduction_7 => 
            next_state <= multiplication_with_reduction_7;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_8;
            end if;
        when multiplication_with_reduction_8 => 
            next_state <= multiplication_with_reduction_8;
            if(penultimate_operation = '1') then
                if(operands_size = "001") then
                    next_state <= multiplication_with_reduction_9;
                else
                    next_state <= multiplication_with_reduction_16;
                end if;
            end if;
        when multiplication_with_reduction_9 => 
            next_state <= multiplication_with_reduction_9;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_10;
            end if;
        when multiplication_with_reduction_10 => 
            next_state <= multiplication_with_reduction_10;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_11;
            end if;
        when multiplication_with_reduction_11 => 
            next_state <= multiplication_with_reduction_11;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_12;
            end if;
        when multiplication_with_reduction_12 => 
            next_state <= multiplication_with_reduction_12;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_13;
            end if;
        when multiplication_with_reduction_13 => 
            next_state <= multiplication_with_reduction_13;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_14;
            end if;
        when multiplication_with_reduction_14 => 
            next_state <= multiplication_with_reduction_14;
            if(penultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when multiplication_with_reduction_16 => 
            next_state <= multiplication_with_reduction_16;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_17;
            end if;
        when multiplication_with_reduction_17 => 
            next_state <= multiplication_with_reduction_17;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_18;
            end if;
        when multiplication_with_reduction_18 => 
            next_state <= multiplication_with_reduction_18;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_19;
            end if;
        when multiplication_with_reduction_19 => 
            next_state <= multiplication_with_reduction_19;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_20;
            end if;
        when multiplication_with_reduction_20 => 
            next_state <= multiplication_with_reduction_20;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_21;
            end if;
        when multiplication_with_reduction_21 => 
            next_state <= multiplication_with_reduction_21;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_22;
            end if;
        when multiplication_with_reduction_22 => 
            next_state <= multiplication_with_reduction_22;
            if(penultimate_operation = '1') then
                if(operands_size = "010") then
                    next_state <= multiplication_with_reduction_23;
                else
                    next_state <= multiplication_with_reduction_34;
                end if;
            end if;
        when multiplication_with_reduction_23 => 
            next_state <= multiplication_with_reduction_23;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_24;
            end if;
        when multiplication_with_reduction_24 => 
            next_state <= multiplication_with_reduction_24;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_25;
            end if;
        when multiplication_with_reduction_25 => 
            next_state <= multiplication_with_reduction_25;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_26;
            end if;
        when multiplication_with_reduction_26 => 
            next_state <= multiplication_with_reduction_26;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_27;
            end if;
        when multiplication_with_reduction_27 => 
            next_state <= multiplication_with_reduction_27;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_28;
            end if;
        when multiplication_with_reduction_28 => 
            next_state <= multiplication_with_reduction_28;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_29;
            end if;
        when multiplication_with_reduction_29 => 
            next_state <= multiplication_with_reduction_29;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_30;
            end if;
        when multiplication_with_reduction_30 => 
            next_state <= multiplication_with_reduction_30;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_31;
            end if;
        when multiplication_with_reduction_31 => 
            next_state <= multiplication_with_reduction_31;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_32;
            end if;
        when multiplication_with_reduction_32 => 
            next_state <= multiplication_with_reduction_32;
            if(penultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when multiplication_with_reduction_34 => 
            next_state <= multiplication_with_reduction_34;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_35;
            end if;
        when multiplication_with_reduction_35 => 
            next_state <= multiplication_with_reduction_35;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_36;
            end if;
        when multiplication_with_reduction_36 => 
            next_state <= multiplication_with_reduction_36;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_37;
            end if;
        when multiplication_with_reduction_37 => 
            next_state <= multiplication_with_reduction_37;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_38;
            end if;
        when multiplication_with_reduction_38 => 
            next_state <= multiplication_with_reduction_38;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_39;
            end if;
        when multiplication_with_reduction_39 => 
            next_state <= multiplication_with_reduction_39;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_40;
            end if;
        when multiplication_with_reduction_40 => 
            next_state <= multiplication_with_reduction_40;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_41;
            end if;
        when multiplication_with_reduction_41 => 
            next_state <= multiplication_with_reduction_41;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_42;
            end if;
        when multiplication_with_reduction_42 => 
            next_state <= multiplication_with_reduction_42;
            if(penultimate_operation = '1') then
                if(operands_size = "011") then
                    next_state <= multiplication_with_reduction_43;
                else
                    next_state <= multiplication_with_reduction_60;
                end if;
            end if;
        when multiplication_with_reduction_43 => 
            next_state <= multiplication_with_reduction_43;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_44;
            end if;
        when multiplication_with_reduction_44 => 
            next_state <= multiplication_with_reduction_44;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_45;
            end if;
        when multiplication_with_reduction_45 => 
            next_state <= multiplication_with_reduction_45;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_46;
            end if;
        when multiplication_with_reduction_46 => 
            next_state <= multiplication_with_reduction_46;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_47;
            end if;
        when multiplication_with_reduction_47 => 
            next_state <= multiplication_with_reduction_47;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_48;
            end if;
        when multiplication_with_reduction_48 => 
            next_state <= multiplication_with_reduction_48;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_49;
            end if;
        when multiplication_with_reduction_49 => 
            next_state <= multiplication_with_reduction_49;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_50;
            end if;
        when multiplication_with_reduction_50 => 
            next_state <= multiplication_with_reduction_50;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_51;
            end if;
        when multiplication_with_reduction_51 => 
            next_state <= multiplication_with_reduction_51;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_52;
            end if;
        when multiplication_with_reduction_52 => 
            next_state <= multiplication_with_reduction_52;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_53;
            end if;
        when multiplication_with_reduction_53 => 
            next_state <= multiplication_with_reduction_53;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_54;
            end if;
        when multiplication_with_reduction_54 => 
            next_state <= multiplication_with_reduction_54;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_55;
            end if;
        when multiplication_with_reduction_55 => 
            next_state <= multiplication_with_reduction_55;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_56;
            end if;
        when multiplication_with_reduction_56 => 
            next_state <= multiplication_with_reduction_56;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_57;
            end if;
        when multiplication_with_reduction_57 => 
            next_state <= multiplication_with_reduction_57;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_58;
            end if;
        when multiplication_with_reduction_58 => 
            next_state <= multiplication_with_reduction_58;
            if(penultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when multiplication_with_reduction_60 => 
            next_state <= multiplication_with_reduction_60;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_61;
            end if;
        when multiplication_with_reduction_61 => 
            next_state <= multiplication_with_reduction_61;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_62;
            end if;
        when multiplication_with_reduction_62 => 
            next_state <= multiplication_with_reduction_62;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_63;
            end if;
        when multiplication_with_reduction_63 => 
            next_state <= multiplication_with_reduction_63;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_64;
            end if;
        when multiplication_with_reduction_64 => 
            next_state <= multiplication_with_reduction_64;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_65;
            end if;
        when multiplication_with_reduction_65 => 
            next_state <= multiplication_with_reduction_65;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_66;
            end if;
        when multiplication_with_reduction_66 => 
            next_state <= multiplication_with_reduction_66;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_67;
            end if;
        when multiplication_with_reduction_67 => 
            next_state <= multiplication_with_reduction_67;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_68;
            end if;
        when multiplication_with_reduction_68 => 
            next_state <= multiplication_with_reduction_68;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_69;
            end if;
        when multiplication_with_reduction_69 => 
            next_state <= multiplication_with_reduction_69;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_70;
            end if;
        when multiplication_with_reduction_70 => 
            next_state <= multiplication_with_reduction_70;
            if(penultimate_operation = '1') then
                if(operands_size = "100") then
                    next_state <= multiplication_with_reduction_71;
                else
                    next_state <= multiplication_with_reduction_96;
                end if;
            end if;
        when multiplication_with_reduction_71 => 
            next_state <= multiplication_with_reduction_71;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_72;
            end if;
        when multiplication_with_reduction_72 => 
            next_state <= multiplication_with_reduction_72;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_73;
            end if;
        when multiplication_with_reduction_73 => 
            next_state <= multiplication_with_reduction_73;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_74;
            end if;
        when multiplication_with_reduction_74 => 
            next_state <= multiplication_with_reduction_74;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_75;
            end if;
        when multiplication_with_reduction_75 => 
            next_state <= multiplication_with_reduction_75;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_76;
            end if;
        when multiplication_with_reduction_76 => 
            next_state <= multiplication_with_reduction_76;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_77;
            end if;
        when multiplication_with_reduction_77 => 
            next_state <= multiplication_with_reduction_77;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_78;
            end if;
        when multiplication_with_reduction_78 => 
            next_state <= multiplication_with_reduction_78;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_79;
            end if;
        when multiplication_with_reduction_79 => 
            next_state <= multiplication_with_reduction_79;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_80;
            end if;
        when multiplication_with_reduction_80 => 
            next_state <= multiplication_with_reduction_80;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_81;
            end if;
        when multiplication_with_reduction_81 => 
            next_state <= multiplication_with_reduction_81;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_82;
            end if;
        when multiplication_with_reduction_82 => 
            next_state <= multiplication_with_reduction_82;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_83;
            end if;
        when multiplication_with_reduction_83 => 
            next_state <= multiplication_with_reduction_83;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_84;
            end if;
        when multiplication_with_reduction_84 => 
            next_state <= multiplication_with_reduction_84;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_85;
            end if;
        when multiplication_with_reduction_85 => 
            next_state <= multiplication_with_reduction_85;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_86;
            end if;
        when multiplication_with_reduction_86 => 
            next_state <= multiplication_with_reduction_86;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_87;
            end if;
        when multiplication_with_reduction_87 => 
            next_state <= multiplication_with_reduction_87;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_88;
            end if;
        when multiplication_with_reduction_88 => 
            next_state <= multiplication_with_reduction_88;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_89;
            end if;
        when multiplication_with_reduction_89 => 
            next_state <= multiplication_with_reduction_89;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_90;
            end if;
        when multiplication_with_reduction_90 => 
            next_state <= multiplication_with_reduction_90;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_91;
            end if;
        when multiplication_with_reduction_91 => 
            next_state <= multiplication_with_reduction_91;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_92;
            end if;
        when multiplication_with_reduction_92 => 
            next_state <= multiplication_with_reduction_92;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_93;
            end if;
        when multiplication_with_reduction_93 => 
            next_state <= multiplication_with_reduction_93;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_94;
            end if;
        when multiplication_with_reduction_94 => 
            next_state <= multiplication_with_reduction_94;
            if(penultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when multiplication_with_reduction_96 => 
            next_state <= multiplication_with_reduction_96;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_97;
            end if;
        when multiplication_with_reduction_97 => 
            next_state <= multiplication_with_reduction_97;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_98;
            end if;
        when multiplication_with_reduction_98 => 
            next_state <= multiplication_with_reduction_98;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_99;
            end if;
        when multiplication_with_reduction_99 => 
            next_state <= multiplication_with_reduction_99;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_100;
            end if;
        when multiplication_with_reduction_100 => 
            next_state <= multiplication_with_reduction_100;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_101;
            end if;
        when multiplication_with_reduction_101 => 
            next_state <= multiplication_with_reduction_101;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_102;
            end if;
        when multiplication_with_reduction_102 => 
            next_state <= multiplication_with_reduction_102;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_103;
            end if;
        when multiplication_with_reduction_103 => 
            next_state <= multiplication_with_reduction_103;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_104;
            end if;
        when multiplication_with_reduction_104 => 
            next_state <= multiplication_with_reduction_104;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_105;
            end if;
        when multiplication_with_reduction_105 => 
            next_state <= multiplication_with_reduction_105;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_106;
            end if;
        when multiplication_with_reduction_106 => 
            next_state <= multiplication_with_reduction_106;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_107;
            end if;
        when multiplication_with_reduction_107 => 
            next_state <= multiplication_with_reduction_107;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_108;
            end if;
        when multiplication_with_reduction_108 => 
            next_state <= multiplication_with_reduction_108;
            if(penultimate_operation = '1') then
                if(operands_size = "101") then
                    next_state <= multiplication_with_reduction_109;
                else
                    next_state <= multiplication_with_reduction_144;
                end if;
            end if;
        when multiplication_with_reduction_109 => 
            next_state <= multiplication_with_reduction_109;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_110;
            end if;
        when multiplication_with_reduction_110 => 
            next_state <= multiplication_with_reduction_110;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_111;
            end if;
        when multiplication_with_reduction_111 => 
            next_state <= multiplication_with_reduction_111;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_112;
            end if;
        when multiplication_with_reduction_112 => 
            next_state <= multiplication_with_reduction_112;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_113;
            end if;
        when multiplication_with_reduction_113 => 
            next_state <= multiplication_with_reduction_113;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_114;
            end if;
        when multiplication_with_reduction_114 => 
            next_state <= multiplication_with_reduction_114;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_115;
            end if;
        when multiplication_with_reduction_115 => 
            next_state <= multiplication_with_reduction_115;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_116;
            end if;
        when multiplication_with_reduction_116 => 
            next_state <= multiplication_with_reduction_116;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_117;
            end if;
        when multiplication_with_reduction_117 => 
            next_state <= multiplication_with_reduction_117;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_118;
            end if;
        when multiplication_with_reduction_118 => 
            next_state <= multiplication_with_reduction_118;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_119;
            end if;
        when multiplication_with_reduction_119 => 
            next_state <= multiplication_with_reduction_119;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_120;
            end if;
        when multiplication_with_reduction_120 => 
            next_state <= multiplication_with_reduction_120;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_121;
            end if;
        when multiplication_with_reduction_121 => 
            next_state <= multiplication_with_reduction_121;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_122;
            end if;
        when multiplication_with_reduction_122 => 
            next_state <= multiplication_with_reduction_122;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_123;
            end if;
        when multiplication_with_reduction_123 => 
            next_state <= multiplication_with_reduction_123;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_124;
            end if;
        when multiplication_with_reduction_124 => 
            next_state <= multiplication_with_reduction_124;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_125;
            end if;
        when multiplication_with_reduction_125 => 
            next_state <= multiplication_with_reduction_125;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_126;
            end if;
        when multiplication_with_reduction_126 => 
            next_state <= multiplication_with_reduction_126;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_127;
            end if;
        when multiplication_with_reduction_127 => 
            next_state <= multiplication_with_reduction_127;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_128;
            end if;
        when multiplication_with_reduction_128 => 
            next_state <= multiplication_with_reduction_128;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_129;
            end if;
        when multiplication_with_reduction_129 => 
            next_state <= multiplication_with_reduction_129;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_130;
            end if;
        when multiplication_with_reduction_130 => 
            next_state <= multiplication_with_reduction_130;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_131;
            end if;
        when multiplication_with_reduction_131 => 
            next_state <= multiplication_with_reduction_131;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_132;
            end if;
        when multiplication_with_reduction_132 => 
            next_state <= multiplication_with_reduction_132;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_133;
            end if;
        when multiplication_with_reduction_133 => 
            next_state <= multiplication_with_reduction_133;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_134;
            end if;
        when multiplication_with_reduction_134 => 
            next_state <= multiplication_with_reduction_134;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_135;
            end if;
        when multiplication_with_reduction_135 => 
            next_state <= multiplication_with_reduction_135;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_136;
            end if;
        when multiplication_with_reduction_136 => 
            next_state <= multiplication_with_reduction_136;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_137;
            end if;
        when multiplication_with_reduction_137 => 
            next_state <= multiplication_with_reduction_137;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_138;
            end if;
        when multiplication_with_reduction_138 => 
            next_state <= multiplication_with_reduction_138;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_139;
            end if;
        when multiplication_with_reduction_139 => 
            next_state <= multiplication_with_reduction_139;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_140;
            end if;
        when multiplication_with_reduction_140 => 
            next_state <= multiplication_with_reduction_140;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_141;
            end if;
        when multiplication_with_reduction_141 => 
            next_state <= multiplication_with_reduction_141;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_142;
            end if;
        when multiplication_with_reduction_142 => 
            next_state <= multiplication_with_reduction_142;
            if(penultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when multiplication_with_reduction_144 => 
            next_state <= multiplication_with_reduction_144;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_145;
            end if;
        when multiplication_with_reduction_145 => 
            next_state <= multiplication_with_reduction_145;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_146;
            end if;
        when multiplication_with_reduction_146 => 
            next_state <= multiplication_with_reduction_146;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_147;
            end if;
        when multiplication_with_reduction_147 => 
            next_state <= multiplication_with_reduction_147;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_148;
            end if;
        when multiplication_with_reduction_148 => 
            next_state <= multiplication_with_reduction_148;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_149;
            end if;
        when multiplication_with_reduction_149 => 
            next_state <= multiplication_with_reduction_149;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_150;
            end if;
        when multiplication_with_reduction_150 => 
            next_state <= multiplication_with_reduction_150;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_151;
            end if;
        when multiplication_with_reduction_151 => 
            next_state <= multiplication_with_reduction_151;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_152;
            end if;
        when multiplication_with_reduction_152 => 
            next_state <= multiplication_with_reduction_152;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_153;
            end if;
        when multiplication_with_reduction_153 => 
            next_state <= multiplication_with_reduction_153;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_154;
            end if;
        when multiplication_with_reduction_154 => 
            next_state <= multiplication_with_reduction_154;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_155;
            end if;
        when multiplication_with_reduction_155 => 
            next_state <= multiplication_with_reduction_155;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_156;
            end if;
        when multiplication_with_reduction_156 => 
            next_state <= multiplication_with_reduction_156;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_157;
            end if;
        when multiplication_with_reduction_157 => 
            next_state <= multiplication_with_reduction_157;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_158;
            end if;
        when multiplication_with_reduction_158 => 
            next_state <= multiplication_with_reduction_158;
            if(penultimate_operation = '1') then
                if(operands_size = "110") then
                    next_state <= multiplication_with_reduction_159;
                else
                    next_state <= multiplication_with_reduction_206;
                end if;
            end if;
        when multiplication_with_reduction_159 => 
            next_state <= multiplication_with_reduction_159;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_160;
            end if;
        when multiplication_with_reduction_160 => 
            next_state <= multiplication_with_reduction_160;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_161;
            end if;
        when multiplication_with_reduction_161 => 
            next_state <= multiplication_with_reduction_161;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_162;
            end if;
        when multiplication_with_reduction_162 => 
            next_state <= multiplication_with_reduction_162;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_163;
            end if;
        when multiplication_with_reduction_163 => 
            next_state <= multiplication_with_reduction_163;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_164;
            end if;
        when multiplication_with_reduction_164 => 
            next_state <= multiplication_with_reduction_164;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_165;
            end if;
        when multiplication_with_reduction_165 => 
            next_state <= multiplication_with_reduction_165;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_166;
            end if;
        when multiplication_with_reduction_166 => 
            next_state <= multiplication_with_reduction_166;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_167;
            end if;
        when multiplication_with_reduction_167 => 
            next_state <= multiplication_with_reduction_167;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_168;
            end if;
        when multiplication_with_reduction_168 => 
            next_state <= multiplication_with_reduction_168;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_169;
            end if;
        when multiplication_with_reduction_169 => 
            next_state <= multiplication_with_reduction_169;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_170;
            end if;
        when multiplication_with_reduction_170 => 
            next_state <= multiplication_with_reduction_170;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_171;
            end if;
        when multiplication_with_reduction_171 => 
            next_state <= multiplication_with_reduction_171;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_172;
            end if;
        when multiplication_with_reduction_172 => 
            next_state <= multiplication_with_reduction_172;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_173;
            end if;
        when multiplication_with_reduction_173 => 
            next_state <= multiplication_with_reduction_173;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_174;
            end if;
        when multiplication_with_reduction_174 => 
            next_state <= multiplication_with_reduction_174;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_175;
            end if;
        when multiplication_with_reduction_175 => 
            next_state <= multiplication_with_reduction_175;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_176;
            end if;
        when multiplication_with_reduction_176 => 
            next_state <= multiplication_with_reduction_176;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_177;
            end if;
        when multiplication_with_reduction_177 => 
            next_state <= multiplication_with_reduction_177;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_178;
            end if;
        when multiplication_with_reduction_178 => 
            next_state <= multiplication_with_reduction_178;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_179;
            end if;
        when multiplication_with_reduction_179 => 
            next_state <= multiplication_with_reduction_179;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_180;
            end if;
        when multiplication_with_reduction_180 => 
            next_state <= multiplication_with_reduction_180;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_181;
            end if;
        when multiplication_with_reduction_181 => 
            next_state <= multiplication_with_reduction_181;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_182;
            end if;
        when multiplication_with_reduction_182 => 
            next_state <= multiplication_with_reduction_182;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_183;
            end if;
        when multiplication_with_reduction_183 => 
            next_state <= multiplication_with_reduction_183;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_184;
            end if;
        when multiplication_with_reduction_184 => 
            next_state <= multiplication_with_reduction_184;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_185;
            end if;
        when multiplication_with_reduction_185 => 
            next_state <= multiplication_with_reduction_185;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_186;
            end if;
        when multiplication_with_reduction_186 => 
            next_state <= multiplication_with_reduction_186;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_187;
            end if;
        when multiplication_with_reduction_187 => 
            next_state <= multiplication_with_reduction_187;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_188;
            end if;
        when multiplication_with_reduction_188 => 
            next_state <= multiplication_with_reduction_188;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_189;
            end if;
        when multiplication_with_reduction_189 => 
            next_state <= multiplication_with_reduction_189;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_190;
            end if;
        when multiplication_with_reduction_190 => 
            next_state <= multiplication_with_reduction_190;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_191;
            end if;
        when multiplication_with_reduction_191 => 
            next_state <= multiplication_with_reduction_191;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_192;
            end if;
        when multiplication_with_reduction_192 => 
            next_state <= multiplication_with_reduction_192;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_193;
            end if;
        when multiplication_with_reduction_193 => 
            next_state <= multiplication_with_reduction_193;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_194;
            end if;
        when multiplication_with_reduction_194 => 
            next_state <= multiplication_with_reduction_194;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_195;
            end if;
        when multiplication_with_reduction_195 => 
            next_state <= multiplication_with_reduction_195;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_196;
            end if;
        when multiplication_with_reduction_196 => 
            next_state <= multiplication_with_reduction_196;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_197;
            end if;
        when multiplication_with_reduction_197 => 
            next_state <= multiplication_with_reduction_197;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_198;
            end if;
        when multiplication_with_reduction_198 => 
            next_state <= multiplication_with_reduction_198;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_199;
            end if;
        when multiplication_with_reduction_199 => 
            next_state <= multiplication_with_reduction_199;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_200;
            end if;
        when multiplication_with_reduction_200 => 
            next_state <= multiplication_with_reduction_200;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_201;
            end if;
        when multiplication_with_reduction_201 => 
            next_state <= multiplication_with_reduction_201;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_202;
            end if;
        when multiplication_with_reduction_202 => 
            next_state <= multiplication_with_reduction_202;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_203;
            end if;
        when multiplication_with_reduction_203 => 
            next_state <= multiplication_with_reduction_203;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_204;
            end if;
        when multiplication_with_reduction_204 => 
            next_state <= multiplication_with_reduction_204;
            if(penultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when multiplication_with_reduction_206 => 
            next_state <= multiplication_with_reduction_206;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_207;
            end if;
        when multiplication_with_reduction_207 => 
            next_state <= multiplication_with_reduction_207;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_208;
            end if;
        when multiplication_with_reduction_208 => 
            next_state <= multiplication_with_reduction_208;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_209;
            end if;
        when multiplication_with_reduction_209 => 
            next_state <= multiplication_with_reduction_209;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_210;
            end if;
        when multiplication_with_reduction_210 => 
            next_state <= multiplication_with_reduction_210;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_211;
            end if;
        when multiplication_with_reduction_211 => 
            next_state <= multiplication_with_reduction_211;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_212;
            end if;
        when multiplication_with_reduction_212 => 
            next_state <= multiplication_with_reduction_212;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_213;
            end if;
        when multiplication_with_reduction_213 => 
            next_state <= multiplication_with_reduction_213;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_214;
            end if;
        when multiplication_with_reduction_214 => 
            next_state <= multiplication_with_reduction_214;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_215;
            end if;
        when multiplication_with_reduction_215 => 
            next_state <= multiplication_with_reduction_215;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_216;
            end if;
        when multiplication_with_reduction_216 => 
            next_state <= multiplication_with_reduction_216;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_217;
            end if;
        when multiplication_with_reduction_217 => 
            next_state <= multiplication_with_reduction_217;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_218;
            end if;
        when multiplication_with_reduction_218 => 
            next_state <= multiplication_with_reduction_218;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_219;
            end if;
        when multiplication_with_reduction_219 => 
            next_state <= multiplication_with_reduction_219;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_220;
            end if;
        when multiplication_with_reduction_220 => 
            next_state <= multiplication_with_reduction_220;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_221;
            end if;
        when multiplication_with_reduction_221 => 
            next_state <= multiplication_with_reduction_221;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_222;
            end if;
        when multiplication_with_reduction_222 => 
            next_state <= multiplication_with_reduction_222;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_223;
            end if;
        when multiplication_with_reduction_223 => 
            next_state <= multiplication_with_reduction_223;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_224;
            end if;
        when multiplication_with_reduction_224 => 
            next_state <= multiplication_with_reduction_224;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_225;
            end if;
        when multiplication_with_reduction_225 => 
            next_state <= multiplication_with_reduction_225;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_226;
            end if;
        when multiplication_with_reduction_226 => 
            next_state <= multiplication_with_reduction_226;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_227;
            end if;
        when multiplication_with_reduction_227 => 
            next_state <= multiplication_with_reduction_227;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_228;
            end if;
        when multiplication_with_reduction_228 => 
            next_state <= multiplication_with_reduction_228;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_229;
            end if;
        when multiplication_with_reduction_229 => 
            next_state <= multiplication_with_reduction_229;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_230;
            end if;
        when multiplication_with_reduction_230 => 
            next_state <= multiplication_with_reduction_230;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_231;
            end if;
        when multiplication_with_reduction_231 => 
            next_state <= multiplication_with_reduction_231;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_232;
            end if;
        when multiplication_with_reduction_232 => 
            next_state <= multiplication_with_reduction_232;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_233;
            end if;
        when multiplication_with_reduction_233 => 
            next_state <= multiplication_with_reduction_233;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_234;
            end if;
        when multiplication_with_reduction_234 => 
            next_state <= multiplication_with_reduction_234;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_235;
            end if;
        when multiplication_with_reduction_235 => 
            next_state <= multiplication_with_reduction_235;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_236;
            end if;
        when multiplication_with_reduction_236 => 
            next_state <= multiplication_with_reduction_236;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_237;
            end if;
        when multiplication_with_reduction_237 => 
            next_state <= multiplication_with_reduction_237;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_238;
            end if;
        when multiplication_with_reduction_238 => 
            next_state <= multiplication_with_reduction_238;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_239;
            end if;
        when multiplication_with_reduction_239 => 
            next_state <= multiplication_with_reduction_239;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_240;
            end if;
        when multiplication_with_reduction_240 => 
            next_state <= multiplication_with_reduction_240;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_241;
            end if;
        when multiplication_with_reduction_241 => 
            next_state <= multiplication_with_reduction_241;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_242;
            end if;
        when multiplication_with_reduction_242 => 
            next_state <= multiplication_with_reduction_242;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_243;
            end if;
        when multiplication_with_reduction_243 => 
            next_state <= multiplication_with_reduction_243;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_244;
            end if;
        when multiplication_with_reduction_244 => 
            next_state <= multiplication_with_reduction_244;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_245;
            end if;
        when multiplication_with_reduction_245 => 
            next_state <= multiplication_with_reduction_245;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_246;
            end if;
        when multiplication_with_reduction_246 => 
            next_state <= multiplication_with_reduction_246;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_247;
            end if;
        when multiplication_with_reduction_247 => 
            next_state <= multiplication_with_reduction_247;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_248;
            end if;
        when multiplication_with_reduction_248 => 
            next_state <= multiplication_with_reduction_248;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_249;
            end if;
        when multiplication_with_reduction_249 => 
            next_state <= multiplication_with_reduction_249;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_250;
            end if;
        when multiplication_with_reduction_250 => 
            next_state <= multiplication_with_reduction_250;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_251;
            end if;
        when multiplication_with_reduction_251 => 
            next_state <= multiplication_with_reduction_251;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_252;
            end if;
        when multiplication_with_reduction_252 => 
            next_state <= multiplication_with_reduction_252;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_253;
            end if;
        when multiplication_with_reduction_253 => 
            next_state <= multiplication_with_reduction_253;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_254;
            end if;
        when multiplication_with_reduction_254 => 
            next_state <= multiplication_with_reduction_254;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_255;
            end if;
        when multiplication_with_reduction_255 => 
            next_state <= multiplication_with_reduction_255;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_256;
            end if;
        when multiplication_with_reduction_256 => 
            next_state <= multiplication_with_reduction_256;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_257;
            end if;
        when multiplication_with_reduction_257 => 
            next_state <= multiplication_with_reduction_257;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_258;
            end if;
        when multiplication_with_reduction_258 => 
            next_state <= multiplication_with_reduction_258;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_259;
            end if;
        when multiplication_with_reduction_259 => 
            next_state <= multiplication_with_reduction_259;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_260;
            end if;
        when multiplication_with_reduction_260 => 
            next_state <= multiplication_with_reduction_260;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_261;
            end if;
        when multiplication_with_reduction_261 => 
            next_state <= multiplication_with_reduction_261;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_262;
            end if;
        when multiplication_with_reduction_262 => 
            next_state <= multiplication_with_reduction_262;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_263;
            end if;
        when multiplication_with_reduction_263 => 
            next_state <= multiplication_with_reduction_263;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_264;
            end if;
        when multiplication_with_reduction_264 => 
            next_state <= multiplication_with_reduction_264;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_265;
            end if;
        when multiplication_with_reduction_265 => 
            next_state <= multiplication_with_reduction_265;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_266;
            end if;
        when multiplication_with_reduction_266 => 
            next_state <= multiplication_with_reduction_266;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_267;
            end if;
        when multiplication_with_reduction_267 => 
            next_state <= multiplication_with_reduction_267;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_268;
            end if;
        when multiplication_with_reduction_268 => 
            next_state <= multiplication_with_reduction_268;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_269;
            end if;
        when multiplication_with_reduction_269 => 
            next_state <= multiplication_with_reduction_269;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_270;
            end if;
        when multiplication_with_reduction_270 => 
            next_state <= multiplication_with_reduction_270;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_271;
            end if;
        when multiplication_with_reduction_271 => 
            next_state <= multiplication_with_reduction_271;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_272;
            end if;
        when multiplication_with_reduction_272 => 
            next_state <= multiplication_with_reduction_272;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_273;
            end if;
        when multiplication_with_reduction_273 => 
            next_state <= multiplication_with_reduction_273;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_274;
            end if;
        when multiplication_with_reduction_274 => 
            next_state <= multiplication_with_reduction_274;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_275;
            end if;
        when multiplication_with_reduction_275 => 
            next_state <= multiplication_with_reduction_275;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_276;
            end if;
        when multiplication_with_reduction_276 => 
            next_state <= multiplication_with_reduction_276;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_277;
            end if;
        when multiplication_with_reduction_277 => 
            next_state <= multiplication_with_reduction_277;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_278;
            end if;
        when multiplication_with_reduction_278 => 
            next_state <= multiplication_with_reduction_278;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_279;
            end if;
        when multiplication_with_reduction_279 => 
            next_state <= multiplication_with_reduction_279;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_280;
            end if;
        when multiplication_with_reduction_280 => 
            next_state <= multiplication_with_reduction_280;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_281;
            end if;
        when multiplication_with_reduction_281 => 
            next_state <= multiplication_with_reduction_281;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_282;
            end if;
        when multiplication_with_reduction_282 => 
            next_state <= multiplication_with_reduction_282;
            if(penultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when multiplication_with_reduction_special_prime_0 => 
            next_state <= multiplication_with_reduction_special_prime_0;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1;
            end if;
        when multiplication_with_reduction_special_prime_1 => 
            next_state <= multiplication_with_reduction_special_prime_1;
            if(penultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when multiplication_with_reduction_special_prime_3 => 
            next_state <= multiplication_with_reduction_special_prime_3;
            if(penultimate_operation = '1') then
                if(operands_size = "001") then
                    next_state <= multiplication_with_reduction_special_prime_4;
                else
                    next_state <= multiplication_with_reduction_special_prime_10;
                end if;
            end if;
        when multiplication_with_reduction_special_prime_4 => 
            next_state <= multiplication_with_reduction_special_prime_4;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_5;
            end if;
        when multiplication_with_reduction_special_prime_5 => 
            next_state <= multiplication_with_reduction_special_prime_5;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_6;
            end if;
        when multiplication_with_reduction_special_prime_6 => 
            next_state <= multiplication_with_reduction_special_prime_6;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_7;
            end if;
        when multiplication_with_reduction_special_prime_7 => 
            next_state <= multiplication_with_reduction_special_prime_7;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_8;
            end if;
        when multiplication_with_reduction_special_prime_8 => 
            next_state <= multiplication_with_reduction_special_prime_8;
            if(penultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when multiplication_with_reduction_special_prime_10 => 
            next_state <= multiplication_with_reduction_special_prime_10;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_11;
            end if;
        when multiplication_with_reduction_special_prime_11 => 
            next_state <= multiplication_with_reduction_special_prime_11;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_12;
            end if;
        when multiplication_with_reduction_special_prime_12 => 
            next_state <= multiplication_with_reduction_special_prime_12;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_13;
            end if;
        when multiplication_with_reduction_special_prime_13 => 
            next_state <= multiplication_with_reduction_special_prime_13;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_14;
            end if;
        when multiplication_with_reduction_special_prime_14 => 
            next_state <= multiplication_with_reduction_special_prime_14;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_15;
            end if;
        when multiplication_with_reduction_special_prime_15 => 
            next_state <= multiplication_with_reduction_special_prime_15;
            if(penultimate_operation = '1') then
                if(operands_size = "010") then
                    next_state <= multiplication_with_reduction_special_prime_16;
                else
                    next_state <= multiplication_with_reduction_special_prime_25;
                end if;
            end if;
        when multiplication_with_reduction_special_prime_16 => 
            next_state <= multiplication_with_reduction_special_prime_16;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_17;
            end if;
        when multiplication_with_reduction_special_prime_17 => 
            next_state <= multiplication_with_reduction_special_prime_17;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_18;
            end if;
        when multiplication_with_reduction_special_prime_18 => 
            next_state <= multiplication_with_reduction_special_prime_18;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_19;
            end if;
        when multiplication_with_reduction_special_prime_19 => 
            next_state <= multiplication_with_reduction_special_prime_19;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_20;
            end if;
        when multiplication_with_reduction_special_prime_20 => 
            next_state <= multiplication_with_reduction_special_prime_20;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_21;
            end if;
        when multiplication_with_reduction_special_prime_21 => 
            next_state <= multiplication_with_reduction_special_prime_21;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_22;
            end if;
        when multiplication_with_reduction_special_prime_22 => 
            next_state <= multiplication_with_reduction_special_prime_22;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_23;
            end if;
        when multiplication_with_reduction_special_prime_23 => 
            next_state <= multiplication_with_reduction_special_prime_23;
            if(penultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when multiplication_with_reduction_special_prime_25 => 
            next_state <= multiplication_with_reduction_special_prime_25;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_26;
            end if;
        when multiplication_with_reduction_special_prime_26 => 
            next_state <= multiplication_with_reduction_special_prime_26;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_27;
            end if;
        when multiplication_with_reduction_special_prime_27 => 
            next_state <= multiplication_with_reduction_special_prime_27;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_28;
            end if;
        when multiplication_with_reduction_special_prime_28 => 
            next_state <= multiplication_with_reduction_special_prime_28;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_29;
            end if;
        when multiplication_with_reduction_special_prime_29 => 
            next_state <= multiplication_with_reduction_special_prime_29;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_30;
            end if;
        when multiplication_with_reduction_special_prime_30 => 
            next_state <= multiplication_with_reduction_special_prime_30;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_31;
            end if;
        when multiplication_with_reduction_special_prime_31 => 
            next_state <= multiplication_with_reduction_special_prime_31;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_32;
            end if;
        when multiplication_with_reduction_special_prime_32 => 
            next_state <= multiplication_with_reduction_special_prime_32;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_33;
            end if;
        when multiplication_with_reduction_special_prime_33 => 
            next_state <= multiplication_with_reduction_special_prime_33;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_34;
            end if;
        when multiplication_with_reduction_special_prime_34 => 
            next_state <= multiplication_with_reduction_special_prime_34;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_35;
            end if;
        when multiplication_with_reduction_special_prime_35 => 
            next_state <= multiplication_with_reduction_special_prime_35;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_36;
            end if;
        when multiplication_with_reduction_special_prime_36 => 
            next_state <= multiplication_with_reduction_special_prime_36;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_37;
            end if;
        when multiplication_with_reduction_special_prime_37 => 
            next_state <= multiplication_with_reduction_special_prime_37;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_38;
            end if;
        when multiplication_with_reduction_special_prime_38 => 
            next_state <= multiplication_with_reduction_special_prime_38;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_39;
            end if;
        when multiplication_with_reduction_special_prime_39 => 
            next_state <= multiplication_with_reduction_special_prime_39;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_40;
            end if;
        when multiplication_with_reduction_special_prime_40 => 
            next_state <= multiplication_with_reduction_special_prime_40;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_41;
            end if;
        when multiplication_with_reduction_special_prime_41 => 
            next_state <= multiplication_with_reduction_special_prime_41;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_42;
            end if;
        when multiplication_with_reduction_special_prime_42 => 
            next_state <= multiplication_with_reduction_special_prime_42;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_43;
            end if;
        when multiplication_with_reduction_special_prime_43 => 
            next_state <= multiplication_with_reduction_special_prime_43;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_44;
            end if;
        when multiplication_with_reduction_special_prime_44 => 
            next_state <= multiplication_with_reduction_special_prime_44;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_45;
            end if;
        when multiplication_with_reduction_special_prime_45 => 
            next_state <= multiplication_with_reduction_special_prime_45;
            if(penultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when multiplication_with_reduction_special_prime_47 => 
            next_state <= multiplication_with_reduction_special_prime_47;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_48;
            end if;
        when multiplication_with_reduction_special_prime_48 => 
            next_state <= multiplication_with_reduction_special_prime_48;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_49;
            end if;
        when multiplication_with_reduction_special_prime_49 => 
            next_state <= multiplication_with_reduction_special_prime_49;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_50;
            end if;
        when multiplication_with_reduction_special_prime_50 => 
            next_state <= multiplication_with_reduction_special_prime_50;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_51;
            end if;
        when multiplication_with_reduction_special_prime_51 => 
            next_state <= multiplication_with_reduction_special_prime_51;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_52;
            end if;
        when multiplication_with_reduction_special_prime_52 => 
            next_state <= multiplication_with_reduction_special_prime_52;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_53;
            end if;
        when multiplication_with_reduction_special_prime_53 => 
            next_state <= multiplication_with_reduction_special_prime_53;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_54;
            end if;
        when multiplication_with_reduction_special_prime_54 => 
            next_state <= multiplication_with_reduction_special_prime_54;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_55;
            end if;
        when multiplication_with_reduction_special_prime_55 => 
            next_state <= multiplication_with_reduction_special_prime_55;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_56;
            end if;
        when multiplication_with_reduction_special_prime_56 => 
            next_state <= multiplication_with_reduction_special_prime_56;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_57;
            end if;
        when multiplication_with_reduction_special_prime_57 => 
            next_state <= multiplication_with_reduction_special_prime_57;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_58;
            end if;
        when multiplication_with_reduction_special_prime_58 => 
            next_state <= multiplication_with_reduction_special_prime_58;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_59;
            end if;
        when multiplication_with_reduction_special_prime_59 => 
            next_state <= multiplication_with_reduction_special_prime_59;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_60;
            end if;
        when multiplication_with_reduction_special_prime_60 => 
            next_state <= multiplication_with_reduction_special_prime_60;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_61;
            end if;
        when multiplication_with_reduction_special_prime_61 => 
            next_state <= multiplication_with_reduction_special_prime_61;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_62;
            end if;
        when multiplication_with_reduction_special_prime_62 => 
            next_state <= multiplication_with_reduction_special_prime_62;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_63;
            end if;
        when multiplication_with_reduction_special_prime_63 => 
            next_state <= multiplication_with_reduction_special_prime_63;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_64;
            end if;
        when multiplication_with_reduction_special_prime_64 => 
            next_state <= multiplication_with_reduction_special_prime_64;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_65;
            end if;
        when multiplication_with_reduction_special_prime_65 => 
            next_state <= multiplication_with_reduction_special_prime_65;
            if(penultimate_operation = '1') then
                if(operands_size = "100") then
                    next_state <= multiplication_with_reduction_special_prime_66;
                else
                    next_state <= multiplication_with_reduction_special_prime_88;
                end if;
            end if;
        when multiplication_with_reduction_special_prime_66 => 
            next_state <= multiplication_with_reduction_special_prime_66;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_67;
            end if;
        when multiplication_with_reduction_special_prime_67 => 
            next_state <= multiplication_with_reduction_special_prime_67;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_68;
            end if;
        when multiplication_with_reduction_special_prime_68 => 
            next_state <= multiplication_with_reduction_special_prime_68;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_69;
            end if;
        when multiplication_with_reduction_special_prime_69 => 
            next_state <= multiplication_with_reduction_special_prime_69;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_70;
            end if;
        when multiplication_with_reduction_special_prime_70 => 
            next_state <= multiplication_with_reduction_special_prime_70;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_71;
            end if;
        when multiplication_with_reduction_special_prime_71 => 
            next_state <= multiplication_with_reduction_special_prime_71;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_72;
            end if;
        when multiplication_with_reduction_special_prime_72 => 
            next_state <= multiplication_with_reduction_special_prime_72;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_73;
            end if;
        when multiplication_with_reduction_special_prime_73 => 
            next_state <= multiplication_with_reduction_special_prime_73;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_74;
            end if;
        when multiplication_with_reduction_special_prime_74 => 
            next_state <= multiplication_with_reduction_special_prime_74;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_75;
            end if;
        when multiplication_with_reduction_special_prime_75 => 
            next_state <= multiplication_with_reduction_special_prime_75;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_76;
            end if;
        when multiplication_with_reduction_special_prime_76 => 
            next_state <= multiplication_with_reduction_special_prime_76;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_77;
            end if;
        when multiplication_with_reduction_special_prime_77 => 
            next_state <= multiplication_with_reduction_special_prime_77;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_78;
            end if;
        when multiplication_with_reduction_special_prime_78 => 
            next_state <= multiplication_with_reduction_special_prime_78;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_79;
            end if;
        when multiplication_with_reduction_special_prime_79 => 
            next_state <= multiplication_with_reduction_special_prime_79;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_80;
            end if;
        when multiplication_with_reduction_special_prime_80 => 
            next_state <= multiplication_with_reduction_special_prime_80;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_81;
            end if;
        when multiplication_with_reduction_special_prime_81 => 
            next_state <= multiplication_with_reduction_special_prime_81;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_82;
            end if;
        when multiplication_with_reduction_special_prime_82 => 
            next_state <= multiplication_with_reduction_special_prime_82;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_83;
            end if;
        when multiplication_with_reduction_special_prime_83 => 
            next_state <= multiplication_with_reduction_special_prime_83;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_84;
            end if;
        when multiplication_with_reduction_special_prime_84 => 
            next_state <= multiplication_with_reduction_special_prime_84;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_85;
            end if;
        when multiplication_with_reduction_special_prime_85 => 
            next_state <= multiplication_with_reduction_special_prime_85;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_86;
            end if;
        when multiplication_with_reduction_special_prime_86 => 
            next_state <= multiplication_with_reduction_special_prime_86;
            if(penultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when multiplication_with_reduction_special_prime_88 => 
            next_state <= multiplication_with_reduction_special_prime_88;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_89;
            end if;
        when multiplication_with_reduction_special_prime_89 => 
            next_state <= multiplication_with_reduction_special_prime_89;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_90;
            end if;
        when multiplication_with_reduction_special_prime_90 => 
            next_state <= multiplication_with_reduction_special_prime_90;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_91;
            end if;
        when multiplication_with_reduction_special_prime_91 => 
            next_state <= multiplication_with_reduction_special_prime_91;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_92;
            end if;
        when multiplication_with_reduction_special_prime_92 => 
            next_state <= multiplication_with_reduction_special_prime_92;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_93;
            end if;
        when multiplication_with_reduction_special_prime_93 => 
            next_state <= multiplication_with_reduction_special_prime_93;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_94;
            end if;
        when multiplication_with_reduction_special_prime_94 => 
            next_state <= multiplication_with_reduction_special_prime_94;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_95;
            end if;
        when multiplication_with_reduction_special_prime_95 => 
            next_state <= multiplication_with_reduction_special_prime_95;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_96;
            end if;
        when multiplication_with_reduction_special_prime_96 => 
            next_state <= multiplication_with_reduction_special_prime_96;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_97;
            end if;
        when multiplication_with_reduction_special_prime_97 => 
            next_state <= multiplication_with_reduction_special_prime_97;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_98;
            end if;
        when multiplication_with_reduction_special_prime_98 => 
            next_state <= multiplication_with_reduction_special_prime_98;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_99;
            end if;
        when multiplication_with_reduction_special_prime_99 => 
            next_state <= multiplication_with_reduction_special_prime_99;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_100;
            end if;
        when multiplication_with_reduction_special_prime_100 => 
            next_state <= multiplication_with_reduction_special_prime_100;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_101;
            end if;
        when multiplication_with_reduction_special_prime_101 => 
            next_state <= multiplication_with_reduction_special_prime_101;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_102;
            end if;
        when multiplication_with_reduction_special_prime_102 => 
            next_state <= multiplication_with_reduction_special_prime_102;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_103;
            end if;
        when multiplication_with_reduction_special_prime_103 => 
            next_state <= multiplication_with_reduction_special_prime_103;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_104;
            end if;
        when multiplication_with_reduction_special_prime_104 => 
            next_state <= multiplication_with_reduction_special_prime_104;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_105;
            end if;
        when multiplication_with_reduction_special_prime_105 => 
            next_state <= multiplication_with_reduction_special_prime_105;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_106;
            end if;
        when multiplication_with_reduction_special_prime_106 => 
            next_state <= multiplication_with_reduction_special_prime_106;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_107;
            end if;
        when multiplication_with_reduction_special_prime_107 => 
            next_state <= multiplication_with_reduction_special_prime_107;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_108;
            end if;
        when multiplication_with_reduction_special_prime_108 => 
            next_state <= multiplication_with_reduction_special_prime_108;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_109;
            end if;
        when multiplication_with_reduction_special_prime_109 => 
            next_state <= multiplication_with_reduction_special_prime_109;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_110;
            end if;
        when multiplication_with_reduction_special_prime_110 => 
            next_state <= multiplication_with_reduction_special_prime_110;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_111;
            end if;
        when multiplication_with_reduction_special_prime_111 => 
            next_state <= multiplication_with_reduction_special_prime_111;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_112;
            end if;
        when multiplication_with_reduction_special_prime_112 => 
            next_state <= multiplication_with_reduction_special_prime_112;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_113;
            end if;
        when multiplication_with_reduction_special_prime_113 => 
            next_state <= multiplication_with_reduction_special_prime_113;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_114;
            end if;
        when multiplication_with_reduction_special_prime_114 => 
            next_state <= multiplication_with_reduction_special_prime_114;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_115;
            end if;
        when multiplication_with_reduction_special_prime_115 => 
            next_state <= multiplication_with_reduction_special_prime_115;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_116;
            end if;
        when multiplication_with_reduction_special_prime_116 => 
            next_state <= multiplication_with_reduction_special_prime_116;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_117;
            end if;
        when multiplication_with_reduction_special_prime_117 => 
            next_state <= multiplication_with_reduction_special_prime_117;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_118;
            end if;
        when multiplication_with_reduction_special_prime_118 => 
            next_state <= multiplication_with_reduction_special_prime_118;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_119;
            end if;
        when multiplication_with_reduction_special_prime_119 => 
            next_state <= multiplication_with_reduction_special_prime_119;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_120;
            end if;
        when multiplication_with_reduction_special_prime_120 => 
            next_state <= multiplication_with_reduction_special_prime_120;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_121;
            end if;
        when multiplication_with_reduction_special_prime_121 => 
            next_state <= multiplication_with_reduction_special_prime_121;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_122;
            end if;
        when multiplication_with_reduction_special_prime_122 => 
            next_state <= multiplication_with_reduction_special_prime_122;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_123;
            end if;
        when multiplication_with_reduction_special_prime_123 => 
            next_state <= multiplication_with_reduction_special_prime_123;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_124;
            end if;
        when multiplication_with_reduction_special_prime_124 => 
            next_state <= multiplication_with_reduction_special_prime_124;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_125;
            end if;
        when multiplication_with_reduction_special_prime_125 => 
            next_state <= multiplication_with_reduction_special_prime_125;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_126;
            end if;
        when multiplication_with_reduction_special_prime_126 => 
            next_state <= multiplication_with_reduction_special_prime_126;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_127;
            end if;
        when multiplication_with_reduction_special_prime_127 => 
            next_state <= multiplication_with_reduction_special_prime_127;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_128;
            end if;
        when multiplication_with_reduction_special_prime_128 => 
            next_state <= multiplication_with_reduction_special_prime_128;
            if(penultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when multiplication_with_reduction_special_prime_130 =>
            next_state <= multiplication_with_reduction_special_prime_130;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_131;
            end if;
        when multiplication_with_reduction_special_prime_131 =>
            next_state <= multiplication_with_reduction_special_prime_131;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_132;
            end if;
        when multiplication_with_reduction_special_prime_132 =>
            next_state <= multiplication_with_reduction_special_prime_132;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_133;
            end if;
        when multiplication_with_reduction_special_prime_133 =>
            next_state <= multiplication_with_reduction_special_prime_133;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_134;
            end if;
        when multiplication_with_reduction_special_prime_134 =>
            next_state <= multiplication_with_reduction_special_prime_134;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_135;
            end if;
        when multiplication_with_reduction_special_prime_135 =>
            next_state <= multiplication_with_reduction_special_prime_135;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_136;
            end if;
        when multiplication_with_reduction_special_prime_136 =>
            next_state <= multiplication_with_reduction_special_prime_136;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_137;
            end if;
        when multiplication_with_reduction_special_prime_137 =>
            next_state <= multiplication_with_reduction_special_prime_137;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_138;
            end if;
        when multiplication_with_reduction_special_prime_138 =>
            next_state <= multiplication_with_reduction_special_prime_138;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_139;
            end if;
        when multiplication_with_reduction_special_prime_139 =>
            next_state <= multiplication_with_reduction_special_prime_139;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_140;
            end if;
        when multiplication_with_reduction_special_prime_140 =>
            next_state <= multiplication_with_reduction_special_prime_140;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_141;
            end if;
        when multiplication_with_reduction_special_prime_141 =>
            next_state <= multiplication_with_reduction_special_prime_141;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_142;
            end if;
        when multiplication_with_reduction_special_prime_142 =>
            next_state <= multiplication_with_reduction_special_prime_142;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_143;
            end if;
        when multiplication_with_reduction_special_prime_143 =>
            next_state <= multiplication_with_reduction_special_prime_143;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_144;
            end if;
        when multiplication_with_reduction_special_prime_144 =>
            next_state <= multiplication_with_reduction_special_prime_144;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_145;
            end if;
        when multiplication_with_reduction_special_prime_145 =>
            next_state <= multiplication_with_reduction_special_prime_145;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_146;
            end if;
        when multiplication_with_reduction_special_prime_146 =>
            next_state <= multiplication_with_reduction_special_prime_146;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_147;
            end if;
        when multiplication_with_reduction_special_prime_147 =>
            next_state <= multiplication_with_reduction_special_prime_147;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_148;
            end if;
        when multiplication_with_reduction_special_prime_148 =>
            next_state <= multiplication_with_reduction_special_prime_148;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_149;
            end if;
        when multiplication_with_reduction_special_prime_149 =>
            next_state <= multiplication_with_reduction_special_prime_149;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_150;
            end if;
        when multiplication_with_reduction_special_prime_150 =>
            next_state <= multiplication_with_reduction_special_prime_150;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_151;
            end if;
        when multiplication_with_reduction_special_prime_151 =>
            next_state <= multiplication_with_reduction_special_prime_151;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_152;
            end if;
        when multiplication_with_reduction_special_prime_152 =>
            next_state <= multiplication_with_reduction_special_prime_152;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_153;
            end if;
        when multiplication_with_reduction_special_prime_153 =>
            next_state <= multiplication_with_reduction_special_prime_153;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_154;
            end if;
        when multiplication_with_reduction_special_prime_154 =>
            next_state <= multiplication_with_reduction_special_prime_154;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_155;
            end if;
        when multiplication_with_reduction_special_prime_155 =>
            next_state <= multiplication_with_reduction_special_prime_155;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_156;
            end if;
        when multiplication_with_reduction_special_prime_156 =>
            next_state <= multiplication_with_reduction_special_prime_156;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_157;
            end if;
        when multiplication_with_reduction_special_prime_157 =>
            next_state <= multiplication_with_reduction_special_prime_157;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_158;
            end if;
        when multiplication_with_reduction_special_prime_158 =>
            next_state <= multiplication_with_reduction_special_prime_158;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_159;
            end if;
        when multiplication_with_reduction_special_prime_159 =>
            next_state <= multiplication_with_reduction_special_prime_159;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_160;
            end if;
        when multiplication_with_reduction_special_prime_160 =>
            next_state <= multiplication_with_reduction_special_prime_160;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_161;
            end if;
        when multiplication_with_reduction_special_prime_161 =>
            next_state <= multiplication_with_reduction_special_prime_161;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_162;
            end if;
        when multiplication_with_reduction_special_prime_162 =>
            next_state <= multiplication_with_reduction_special_prime_162;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_163;
            end if;
        when multiplication_with_reduction_special_prime_163 =>
            next_state <= multiplication_with_reduction_special_prime_163;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_164;
            end if;
        when multiplication_with_reduction_special_prime_164 =>
            next_state <= multiplication_with_reduction_special_prime_164;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_165;
            end if;
        when multiplication_with_reduction_special_prime_165 => 
            next_state <= multiplication_with_reduction_special_prime_165;
            if(penultimate_operation = '1') then
                if(operands_size = "110") then
                    next_state <= multiplication_with_reduction_special_prime_166;
                else
                    next_state <= multiplication_with_reduction_special_prime_208;
                end if;
                
            end if;
        when multiplication_with_reduction_special_prime_166 => 
            next_state <= multiplication_with_reduction_special_prime_166;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_167;
            end if;
        when multiplication_with_reduction_special_prime_167 => 
            next_state <= multiplication_with_reduction_special_prime_167;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_168;
            end if;
        when multiplication_with_reduction_special_prime_168 => 
            next_state <= multiplication_with_reduction_special_prime_168;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_169;
            end if;
        when multiplication_with_reduction_special_prime_169 => 
            next_state <= multiplication_with_reduction_special_prime_169;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_170;
            end if;
        when multiplication_with_reduction_special_prime_170 => 
            next_state <= multiplication_with_reduction_special_prime_170;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_171;
            end if;
        when multiplication_with_reduction_special_prime_171 => 
            next_state <= multiplication_with_reduction_special_prime_171;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_172;
            end if;
        when multiplication_with_reduction_special_prime_172 => 
            next_state <= multiplication_with_reduction_special_prime_172;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_173;
            end if;
        when multiplication_with_reduction_special_prime_173 => 
            next_state <= multiplication_with_reduction_special_prime_173;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_174;
            end if;
        when multiplication_with_reduction_special_prime_174 => 
            next_state <= multiplication_with_reduction_special_prime_174;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_175;
            end if;
        when multiplication_with_reduction_special_prime_175 => 
            next_state <= multiplication_with_reduction_special_prime_175;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_176;
            end if;
        when multiplication_with_reduction_special_prime_176 => 
            next_state <= multiplication_with_reduction_special_prime_176;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_177;
            end if;
        when multiplication_with_reduction_special_prime_177 => 
            next_state <= multiplication_with_reduction_special_prime_177;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_178;
            end if;
        when multiplication_with_reduction_special_prime_178 => 
            next_state <= multiplication_with_reduction_special_prime_178;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_179;
            end if;
        when multiplication_with_reduction_special_prime_179 => 
            next_state <= multiplication_with_reduction_special_prime_179;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_180;
            end if;
        when multiplication_with_reduction_special_prime_180 => 
            next_state <= multiplication_with_reduction_special_prime_180;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_181;
            end if;
        when multiplication_with_reduction_special_prime_181 => 
            next_state <= multiplication_with_reduction_special_prime_181;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_182;
            end if;
        when multiplication_with_reduction_special_prime_182 => 
            next_state <= multiplication_with_reduction_special_prime_182;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_183;
            end if;
        when multiplication_with_reduction_special_prime_183 => 
            next_state <= multiplication_with_reduction_special_prime_183;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_184;
            end if;
        when multiplication_with_reduction_special_prime_184 => 
            next_state <= multiplication_with_reduction_special_prime_184;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_185;
            end if;
        when multiplication_with_reduction_special_prime_185 => 
            next_state <= multiplication_with_reduction_special_prime_185;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_186;
            end if;
        when multiplication_with_reduction_special_prime_186 => 
            next_state <= multiplication_with_reduction_special_prime_186;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_187;
            end if;
        when multiplication_with_reduction_special_prime_187 => 
            next_state <= multiplication_with_reduction_special_prime_187;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_188;
            end if;
        when multiplication_with_reduction_special_prime_188 => 
            next_state <= multiplication_with_reduction_special_prime_188;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_189;
            end if;
        when multiplication_with_reduction_special_prime_189 => 
            next_state <= multiplication_with_reduction_special_prime_189;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_190;
            end if;
        when multiplication_with_reduction_special_prime_190 => 
            next_state <= multiplication_with_reduction_special_prime_190;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_191;
            end if;
        when multiplication_with_reduction_special_prime_191 => 
            next_state <= multiplication_with_reduction_special_prime_191;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_192;
            end if;
        when multiplication_with_reduction_special_prime_192 => 
            next_state <= multiplication_with_reduction_special_prime_192;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_193;
            end if;
        when multiplication_with_reduction_special_prime_193 => 
            next_state <= multiplication_with_reduction_special_prime_193;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_194;
            end if;
        when multiplication_with_reduction_special_prime_194 => 
            next_state <= multiplication_with_reduction_special_prime_194;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_195;
            end if;
        when multiplication_with_reduction_special_prime_195 => 
            next_state <= multiplication_with_reduction_special_prime_195;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_196;
            end if;
        when multiplication_with_reduction_special_prime_196 => 
            next_state <= multiplication_with_reduction_special_prime_196;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_197;
            end if;
        when multiplication_with_reduction_special_prime_197 => 
            next_state <= multiplication_with_reduction_special_prime_197;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_198;
            end if;
        when multiplication_with_reduction_special_prime_198 => 
            next_state <= multiplication_with_reduction_special_prime_198;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_199;
            end if;
        when multiplication_with_reduction_special_prime_199 => 
            next_state <= multiplication_with_reduction_special_prime_199;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_200;
            end if;
        when multiplication_with_reduction_special_prime_200 => 
            next_state <= multiplication_with_reduction_special_prime_200;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_201;
            end if;
        when multiplication_with_reduction_special_prime_201 => 
            next_state <= multiplication_with_reduction_special_prime_201;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_202;
            end if;
        when multiplication_with_reduction_special_prime_202 => 
            next_state <= multiplication_with_reduction_special_prime_202;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_203;
            end if;
        when multiplication_with_reduction_special_prime_203 => 
            next_state <= multiplication_with_reduction_special_prime_203;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_204;
            end if;
        when multiplication_with_reduction_special_prime_204 => 
            next_state <= multiplication_with_reduction_special_prime_204;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_205;
            end if;
        when multiplication_with_reduction_special_prime_205 => 
            next_state <= multiplication_with_reduction_special_prime_205;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_206;
            end if;
        when multiplication_with_reduction_special_prime_206 => 
            next_state <= multiplication_with_reduction_special_prime_206;
            if(penultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when multiplication_with_reduction_special_prime_208 => 
            next_state <= multiplication_with_reduction_special_prime_208;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_209;
            end if;
        when multiplication_with_reduction_special_prime_209 => 
            next_state <= multiplication_with_reduction_special_prime_209;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_210;
            end if;
        when multiplication_with_reduction_special_prime_210 => 
            next_state <= multiplication_with_reduction_special_prime_210;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_211;
            end if;
        when multiplication_with_reduction_special_prime_211 => 
            next_state <= multiplication_with_reduction_special_prime_211;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_212;
            end if;
        when multiplication_with_reduction_special_prime_212 => 
            next_state <= multiplication_with_reduction_special_prime_212;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_213;
            end if;
        when multiplication_with_reduction_special_prime_213 => 
            next_state <= multiplication_with_reduction_special_prime_213;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_214;
            end if;
        when multiplication_with_reduction_special_prime_214 => 
            next_state <= multiplication_with_reduction_special_prime_214;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_215;
            end if;
        when multiplication_with_reduction_special_prime_215 => 
            next_state <= multiplication_with_reduction_special_prime_215;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_216;
            end if;
        when multiplication_with_reduction_special_prime_216 => 
            next_state <= multiplication_with_reduction_special_prime_216;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_217;
            end if;
        when multiplication_with_reduction_special_prime_217 => 
            next_state <= multiplication_with_reduction_special_prime_217;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_218;
            end if;
        when multiplication_with_reduction_special_prime_218 => 
            next_state <= multiplication_with_reduction_special_prime_218;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_219;
            end if;
        when multiplication_with_reduction_special_prime_219 => 
            next_state <= multiplication_with_reduction_special_prime_219;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_220;
            end if;
        when multiplication_with_reduction_special_prime_220 => 
            next_state <= multiplication_with_reduction_special_prime_220;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_221;
            end if;
        when multiplication_with_reduction_special_prime_221 => 
            next_state <= multiplication_with_reduction_special_prime_221;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_222;
            end if;
        when multiplication_with_reduction_special_prime_222 => 
            next_state <= multiplication_with_reduction_special_prime_222;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_223;
            end if;
        when multiplication_with_reduction_special_prime_223 => 
            next_state <= multiplication_with_reduction_special_prime_223;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_224;
            end if;
        when multiplication_with_reduction_special_prime_224 => 
            next_state <= multiplication_with_reduction_special_prime_224;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_225;
            end if;
        when multiplication_with_reduction_special_prime_225 => 
            next_state <= multiplication_with_reduction_special_prime_225;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_226;
            end if;
        when multiplication_with_reduction_special_prime_226 => 
            next_state <= multiplication_with_reduction_special_prime_226;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_227;
            end if;
        when multiplication_with_reduction_special_prime_227 => 
            next_state <= multiplication_with_reduction_special_prime_227;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_228;
            end if;
        when multiplication_with_reduction_special_prime_228 => 
            next_state <= multiplication_with_reduction_special_prime_228;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_229;
            end if;
        when multiplication_with_reduction_special_prime_229 => 
            next_state <= multiplication_with_reduction_special_prime_229;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_230;
            end if;
        when multiplication_with_reduction_special_prime_230 => 
            next_state <= multiplication_with_reduction_special_prime_230;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_231;
            end if;
        when multiplication_with_reduction_special_prime_231 => 
            next_state <= multiplication_with_reduction_special_prime_231;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_232;
            end if;
        when multiplication_with_reduction_special_prime_232 => 
            next_state <= multiplication_with_reduction_special_prime_232;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_233;
            end if;
        when multiplication_with_reduction_special_prime_233 => 
            next_state <= multiplication_with_reduction_special_prime_233;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_234;
            end if;
        when multiplication_with_reduction_special_prime_234 => 
            next_state <= multiplication_with_reduction_special_prime_234;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_235;
            end if;
        when multiplication_with_reduction_special_prime_235 => 
            next_state <= multiplication_with_reduction_special_prime_235;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_236;
            end if;
        when multiplication_with_reduction_special_prime_236 => 
            next_state <= multiplication_with_reduction_special_prime_236;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_237;
            end if;
        when multiplication_with_reduction_special_prime_237 => 
            next_state <= multiplication_with_reduction_special_prime_237;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_238;
            end if;
        when multiplication_with_reduction_special_prime_238 => 
            next_state <= multiplication_with_reduction_special_prime_238;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_239;
            end if;
        when multiplication_with_reduction_special_prime_239 => 
            next_state <= multiplication_with_reduction_special_prime_239;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_240;
            end if;
        when multiplication_with_reduction_special_prime_240 => 
            next_state <= multiplication_with_reduction_special_prime_240;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_241;
            end if;
        when multiplication_with_reduction_special_prime_241 => 
            next_state <= multiplication_with_reduction_special_prime_241;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_242;
            end if;
        when multiplication_with_reduction_special_prime_242 => 
            next_state <= multiplication_with_reduction_special_prime_242;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_243;
            end if;
        when multiplication_with_reduction_special_prime_243 => 
            next_state <= multiplication_with_reduction_special_prime_243;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_244;
            end if;
        when multiplication_with_reduction_special_prime_244 => 
            next_state <= multiplication_with_reduction_special_prime_244;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_245;
            end if;
        when multiplication_with_reduction_special_prime_245 => 
            next_state <= multiplication_with_reduction_special_prime_245;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_246;
            end if;
        when multiplication_with_reduction_special_prime_246 => 
            next_state <= multiplication_with_reduction_special_prime_246;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_247;
            end if;
        when multiplication_with_reduction_special_prime_247 => 
            next_state <= multiplication_with_reduction_special_prime_247;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_248;
            end if;
        when multiplication_with_reduction_special_prime_248 => 
            next_state <= multiplication_with_reduction_special_prime_248;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_249;
            end if;
        when multiplication_with_reduction_special_prime_249 => 
            next_state <= multiplication_with_reduction_special_prime_249;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_250;
            end if;
        when multiplication_with_reduction_special_prime_250 => 
            next_state <= multiplication_with_reduction_special_prime_250;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_251;
            end if;
        when multiplication_with_reduction_special_prime_251 => 
            next_state <= multiplication_with_reduction_special_prime_251;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_252;
            end if;
        when multiplication_with_reduction_special_prime_252 => 
            next_state <= multiplication_with_reduction_special_prime_252;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_253;
            end if;
        when multiplication_with_reduction_special_prime_253 => 
            next_state <= multiplication_with_reduction_special_prime_253;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_254;
            end if;
        when multiplication_with_reduction_special_prime_254 => 
            next_state <= multiplication_with_reduction_special_prime_254;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_255;
            end if;
        when multiplication_with_reduction_special_prime_255 => 
            next_state <= multiplication_with_reduction_special_prime_255;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_256;
            end if;
        when multiplication_with_reduction_special_prime_256 => 
            next_state <= multiplication_with_reduction_special_prime_256;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_257;
            end if;
        when multiplication_with_reduction_special_prime_257 => 
            next_state <= multiplication_with_reduction_special_prime_257;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_258;
            end if;
        when multiplication_with_reduction_special_prime_258 => 
            next_state <= multiplication_with_reduction_special_prime_258;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_259;
            end if;
        when multiplication_with_reduction_special_prime_259 => 
            next_state <= multiplication_with_reduction_special_prime_259;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_260;
            end if;
        when multiplication_with_reduction_special_prime_260 => 
            next_state <= multiplication_with_reduction_special_prime_260;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_261;
            end if;
        when multiplication_with_reduction_special_prime_261 => 
            next_state <= multiplication_with_reduction_special_prime_261;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_262;
            end if;
        when multiplication_with_reduction_special_prime_262 => 
            next_state <= multiplication_with_reduction_special_prime_262;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_263;
            end if;
        when multiplication_with_reduction_special_prime_263 => 
            next_state <= multiplication_with_reduction_special_prime_263;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_264;
            end if;
        when multiplication_with_reduction_special_prime_264 => 
            next_state <= multiplication_with_reduction_special_prime_264;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_265;
            end if;
        when multiplication_with_reduction_special_prime_265 => 
            next_state <= multiplication_with_reduction_special_prime_265;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_266;
            end if;
        when multiplication_with_reduction_special_prime_266 => 
            next_state <= multiplication_with_reduction_special_prime_266;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_267;
            end if;
        when multiplication_with_reduction_special_prime_267 => 
            next_state <= multiplication_with_reduction_special_prime_267;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_268;
            end if;
        when multiplication_with_reduction_special_prime_268 => 
            next_state <= multiplication_with_reduction_special_prime_268;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_269;
            end if;
        when multiplication_with_reduction_special_prime_269 => 
            next_state <= multiplication_with_reduction_special_prime_269;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_270;
            end if;
        when multiplication_with_reduction_special_prime_270 => 
            next_state <= multiplication_with_reduction_special_prime_270;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_271;
            end if;
        when multiplication_with_reduction_special_prime_271 => 
            next_state <= multiplication_with_reduction_special_prime_271;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_272;
            end if;
        when multiplication_with_reduction_special_prime_272 => 
            next_state <= multiplication_with_reduction_special_prime_272;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_273;
            end if;
        when multiplication_with_reduction_special_prime_273 => 
            next_state <= multiplication_with_reduction_special_prime_273;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_274;
            end if;
        when multiplication_with_reduction_special_prime_274 => 
            next_state <= multiplication_with_reduction_special_prime_274;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_275;
            end if;
        when multiplication_with_reduction_special_prime_275 => 
            next_state <= multiplication_with_reduction_special_prime_275;
            if(penultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when square_with_reduction_0 => 
            next_state <= square_with_reduction_0;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_1;
            end if;
        when square_with_reduction_1 => 
            next_state <= square_with_reduction_1;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_2;
            end if;
        when square_with_reduction_2 => 
            next_state <= square_with_reduction_2;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_3;
            end if;
        when square_with_reduction_3 => 
            next_state <= square_with_reduction_3;
            if(penultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when square_with_reduction_5 => 
            next_state <= square_with_reduction_5;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_6;
            end if;
        when square_with_reduction_6 => 
            next_state <= square_with_reduction_6;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_7;
            end if;
        when square_with_reduction_7 => 
            next_state <= square_with_reduction_7;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_8;
            end if;
        when square_with_reduction_8 => 
            next_state <= square_with_reduction_8;
            if(penultimate_operation = '1') then
                if(operands_size = "001") then
                    next_state <= square_with_reduction_9;
                else
                    next_state <= square_with_reduction_15;
                end if;
            end if;
        when square_with_reduction_9 => 
            next_state <= square_with_reduction_9;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_10;
            end if;
        when square_with_reduction_10 => 
            next_state <= square_with_reduction_10;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_11;
            end if;
        when square_with_reduction_11 => 
            next_state <= square_with_reduction_11;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_12;
            end if;
        when square_with_reduction_12 => 
            next_state <= square_with_reduction_12;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_13;
            end if;
        when square_with_reduction_13 => 
            next_state <= square_with_reduction_13;
            if(penultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when square_with_reduction_15 => 
            next_state <= square_with_reduction_15;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_16;
            end if;
        when square_with_reduction_16 => 
            next_state <= square_with_reduction_16;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_17;
            end if;
        when square_with_reduction_17 => 
            next_state <= square_with_reduction_17;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_18;
            end if;
        when square_with_reduction_18 => 
            next_state <= square_with_reduction_18;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_19;
            end if;
        when square_with_reduction_19 => 
            next_state <= square_with_reduction_19;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_20;
            end if;
        when square_with_reduction_20 => 
            next_state <= square_with_reduction_20;
            if(penultimate_operation = '1') then
                if(operands_size = "010") then
                    next_state <= square_with_reduction_21;
                else
                    next_state <= square_with_reduction_30;
                end if;
            end if;
        when square_with_reduction_21 => 
            next_state <= square_with_reduction_21;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_22;
            end if;
        when square_with_reduction_22 => 
            next_state <= square_with_reduction_22;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_23;
            end if;
        when square_with_reduction_23 => 
            next_state <= square_with_reduction_23;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_24;
            end if;
        when square_with_reduction_24 => 
            next_state <= square_with_reduction_24;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_25;
            end if;
        when square_with_reduction_25 => 
            next_state <= square_with_reduction_25;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_26;
            end if;
        when square_with_reduction_26 => 
            next_state <= square_with_reduction_26;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_27;
            end if;
        when square_with_reduction_27 => 
            next_state <= square_with_reduction_27;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_28;
            end if;
        when square_with_reduction_28 => 
            next_state <= square_with_reduction_28;
            if(penultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when square_with_reduction_30 => 
            next_state <= square_with_reduction_30;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_31;
            end if;
        when square_with_reduction_31 => 
            next_state <= square_with_reduction_31;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_32;
            end if;
        when square_with_reduction_32 => 
            next_state <= square_with_reduction_32;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_33;
            end if;
        when square_with_reduction_33 => 
            next_state <= square_with_reduction_33;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_34;
            end if;
        when square_with_reduction_34 => 
            next_state <= square_with_reduction_34;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_35;
            end if;
        when square_with_reduction_35 => 
            next_state <= square_with_reduction_35;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_36;
            end if;
        when square_with_reduction_36 => 
            next_state <= square_with_reduction_36;
            if(penultimate_operation = '1') then
                if(operands_size = "011") then
                    next_state <= square_with_reduction_37;
                else
                    next_state <= square_with_reduction_51;
                end if;
            end if;
        when square_with_reduction_37 => 
            next_state <= square_with_reduction_37;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_38;
            end if;
        when square_with_reduction_38 => 
            next_state <= square_with_reduction_38;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_39;
            end if;
        when square_with_reduction_39 => 
            next_state <= square_with_reduction_39;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_40;
            end if;
        when square_with_reduction_40 => 
            next_state <= square_with_reduction_40;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_41;
            end if;
        when square_with_reduction_41 => 
            next_state <= square_with_reduction_41;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_42;
            end if;
        when square_with_reduction_42 => 
            next_state <= square_with_reduction_42;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_43;
            end if;
        when square_with_reduction_43 => 
            next_state <= square_with_reduction_43;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_44;
            end if;
        when square_with_reduction_44 => 
            next_state <= square_with_reduction_44;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_45;
            end if;
        when square_with_reduction_45 => 
            next_state <= square_with_reduction_45;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_46;
            end if;
        when square_with_reduction_46 => 
            next_state <= square_with_reduction_46;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_47;
            end if;
        when square_with_reduction_47 => 
            next_state <= square_with_reduction_47;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_48;
            end if;
        when square_with_reduction_48 => 
            next_state <= square_with_reduction_48;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_49;
            end if;
        when square_with_reduction_49 => 
            next_state <= square_with_reduction_49;
            if(penultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when square_with_reduction_51 => 
            next_state <= square_with_reduction_51;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_52;
            end if;
        when square_with_reduction_52 => 
            next_state <= square_with_reduction_52;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_53;
            end if;
        when square_with_reduction_53 => 
            next_state <= square_with_reduction_53;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_54;
            end if;
        when square_with_reduction_54 => 
            next_state <= square_with_reduction_54;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_55;
            end if;
        when square_with_reduction_55 => 
            next_state <= square_with_reduction_55;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_56;
            end if;
        when square_with_reduction_56 => 
            next_state <= square_with_reduction_56;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_57;
            end if;
        when square_with_reduction_57 => 
            next_state <= square_with_reduction_57;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_58;
            end if;
        when square_with_reduction_58 => 
            next_state <= square_with_reduction_58;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_59;
            end if;
        when square_with_reduction_59 => 
            next_state <= square_with_reduction_59;
            if(penultimate_operation = '1') then
                if(operands_size = "100") then
                    next_state <= square_with_reduction_60;
                else
                    next_state <= square_with_reduction_80;
                end if;
            end if;
        when square_with_reduction_60 => 
            next_state <= square_with_reduction_60;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_61;
            end if;
        when square_with_reduction_61 => 
            next_state <= square_with_reduction_61;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_62;
            end if;
        when square_with_reduction_62 => 
            next_state <= square_with_reduction_62;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_63;
            end if;
        when square_with_reduction_63 => 
            next_state <= square_with_reduction_63;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_64;
            end if;
        when square_with_reduction_64 => 
            next_state <= square_with_reduction_64;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_65;
            end if;
        when square_with_reduction_65 => 
            next_state <= square_with_reduction_65;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_66;
            end if;
        when square_with_reduction_66 => 
            next_state <= square_with_reduction_66;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_67;
            end if;
        when square_with_reduction_67 => 
            next_state <= square_with_reduction_67;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_68;
            end if;
        when square_with_reduction_68 => 
            next_state <= square_with_reduction_68;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_69;
            end if;
        when square_with_reduction_69 => 
            next_state <= square_with_reduction_69;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_70;
            end if;
        when square_with_reduction_70 => 
            next_state <= square_with_reduction_70;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_71;
            end if;
        when square_with_reduction_71 => 
            next_state <= square_with_reduction_71;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_72;
            end if;
        when square_with_reduction_72 => 
            next_state <= square_with_reduction_72;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_73;
            end if;
        when square_with_reduction_73 => 
            next_state <= square_with_reduction_73;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_74;
            end if;
        when square_with_reduction_74 => 
            next_state <= square_with_reduction_74;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_75;
            end if;
        when square_with_reduction_75 => 
            next_state <= square_with_reduction_75;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_76;
            end if;
        when square_with_reduction_76 => 
            next_state <= square_with_reduction_76;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_77;
            end if;
        when square_with_reduction_77 => 
            next_state <= square_with_reduction_77;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_78;
            end if;
        when square_with_reduction_78 => 
            next_state <= square_with_reduction_78;
            if(penultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when square_with_reduction_80 => 
            next_state <= square_with_reduction_80;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_81;
            end if;
        when square_with_reduction_81 => 
            next_state <= square_with_reduction_81;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_82;
            end if;
        when square_with_reduction_82 => 
            next_state <= square_with_reduction_82;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_83;
            end if;
        when square_with_reduction_83 => 
            next_state <= square_with_reduction_83;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_84;
            end if;
        when square_with_reduction_84 => 
            next_state <= square_with_reduction_84;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_85;
            end if;
        when square_with_reduction_85 => 
            next_state <= square_with_reduction_85;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_86;
            end if;
        when square_with_reduction_86 => 
            next_state <= square_with_reduction_86;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_87;
            end if;
        when square_with_reduction_87 => 
            next_state <= square_with_reduction_87;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_88;
            end if;
        when square_with_reduction_88 => 
            next_state <= square_with_reduction_88;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_89;
            end if;
        when square_with_reduction_89 => 
            next_state <= square_with_reduction_89;
            if(penultimate_operation = '1') then
                if(operands_size = "101") then
                    next_state <= square_with_reduction_90;
                else
                    next_state <= square_with_reduction_118;
                end if;
            end if;
        when square_with_reduction_90 => 
            next_state <= square_with_reduction_90;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_91;
            end if;
        when square_with_reduction_91 => 
            next_state <= square_with_reduction_91;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_92;
            end if;
        when square_with_reduction_92 => 
            next_state <= square_with_reduction_92;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_93;
            end if;
        when square_with_reduction_93 => 
            next_state <= square_with_reduction_93;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_94;
            end if;
        when square_with_reduction_94 => 
            next_state <= square_with_reduction_94;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_95;
            end if;
        when square_with_reduction_95 => 
            next_state <= square_with_reduction_95;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_96;
            end if;
        when square_with_reduction_96 => 
            next_state <= square_with_reduction_96;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_97;
            end if;
        when square_with_reduction_97 => 
            next_state <= square_with_reduction_97;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_98;
            end if;
        when square_with_reduction_98 => 
            next_state <= square_with_reduction_98;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_99;
            end if;
        when square_with_reduction_99 => 
            next_state <= square_with_reduction_99;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_100;
            end if;
        when square_with_reduction_100 => 
            next_state <= square_with_reduction_100;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_101;
            end if;
        when square_with_reduction_101 => 
            next_state <= square_with_reduction_101;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_102;
            end if;
        when square_with_reduction_102 => 
            next_state <= square_with_reduction_102;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_103;
            end if;
        when square_with_reduction_103 => 
            next_state <= square_with_reduction_103;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_104;
            end if;
        when square_with_reduction_104 => 
            next_state <= square_with_reduction_104;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_105;
            end if;
        when square_with_reduction_105 => 
            next_state <= square_with_reduction_105;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_106;
            end if;
        when square_with_reduction_106 => 
            next_state <= square_with_reduction_106;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_107;
            end if;
        when square_with_reduction_107 => 
            next_state <= square_with_reduction_107;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_108;
            end if;
        when square_with_reduction_108 => 
            next_state <= square_with_reduction_108;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_109;
            end if;
        when square_with_reduction_109 => 
            next_state <= square_with_reduction_109;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_110;
            end if;
        when square_with_reduction_110 => 
            next_state <= square_with_reduction_110;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_111;
            end if;
        when square_with_reduction_111 => 
            next_state <= square_with_reduction_111;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_112;
            end if;
        when square_with_reduction_112 => 
            next_state <= square_with_reduction_112;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_113;
            end if;
        when square_with_reduction_113 => 
            next_state <= square_with_reduction_113;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_114;
            end if;
        when square_with_reduction_114 => 
            next_state <= square_with_reduction_114;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_115;
            end if;
        when square_with_reduction_115 => 
            next_state <= square_with_reduction_115;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_116;
            end if;
        when square_with_reduction_116 => 
            next_state <= square_with_reduction_116;
            if(penultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when square_with_reduction_118 => 
            next_state <= square_with_reduction_118;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_119;
            end if;
        when square_with_reduction_119 => 
            next_state <= square_with_reduction_119;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_120;
            end if;
        when square_with_reduction_120 => 
            next_state <= square_with_reduction_120;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_121;
            end if;
        when square_with_reduction_121 => 
            next_state <= square_with_reduction_121;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_122;
            end if;
        when square_with_reduction_122 => 
            next_state <= square_with_reduction_122;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_123;
            end if;
        when square_with_reduction_123 => 
            next_state <= square_with_reduction_123;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_124;
            end if;
        when square_with_reduction_124 => 
            next_state <= square_with_reduction_124;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_125;
            end if;
        when square_with_reduction_125 => 
            next_state <= square_with_reduction_125;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_126;
            end if;
        when square_with_reduction_126 => 
            next_state <= square_with_reduction_126;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_127;
            end if;
        when square_with_reduction_127 => 
            next_state <= square_with_reduction_127;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_128;
            end if;
        when square_with_reduction_128 => 
            next_state <= square_with_reduction_128;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_129;
            end if;
        when square_with_reduction_129 => 
            next_state <= square_with_reduction_129;
            if(penultimate_operation = '1') then
                if(operands_size = "110") then
                    next_state <= square_with_reduction_130;
                else
                    next_state <= square_with_reduction_167;
                end if;
            end if;
        when square_with_reduction_130 => 
            next_state <= square_with_reduction_130;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_131;
            end if;
        when square_with_reduction_131 => 
            next_state <= square_with_reduction_131;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_132;
            end if;
        when square_with_reduction_132 => 
            next_state <= square_with_reduction_132;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_133;
            end if;
        when square_with_reduction_133 => 
            next_state <= square_with_reduction_133;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_134;
            end if;
        when square_with_reduction_134 => 
            next_state <= square_with_reduction_134;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_135;
            end if;
        when square_with_reduction_135 => 
            next_state <= square_with_reduction_135;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_136;
            end if;
        when square_with_reduction_136 => 
            next_state <= square_with_reduction_136;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_137;
            end if;
        when square_with_reduction_137 => 
            next_state <= square_with_reduction_137;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_138;
            end if;
        when square_with_reduction_138 => 
            next_state <= square_with_reduction_138;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_139;
            end if;
        when square_with_reduction_139 => 
            next_state <= square_with_reduction_139;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_140;
            end if;
        when square_with_reduction_140 => 
            next_state <= square_with_reduction_140;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_141;
            end if;
        when square_with_reduction_141 => 
            next_state <= square_with_reduction_141;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_142;
            end if;
        when square_with_reduction_142 => 
            next_state <= square_with_reduction_142;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_143;
            end if;
        when square_with_reduction_143 => 
            next_state <= square_with_reduction_143;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_144;
            end if;
        when square_with_reduction_144 => 
            next_state <= square_with_reduction_144;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_145;
            end if;
        when square_with_reduction_145 => 
            next_state <= square_with_reduction_145;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_146;
            end if;
        when square_with_reduction_146 => 
            next_state <= square_with_reduction_146;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_147;
            end if;
        when square_with_reduction_147 => 
            next_state <= square_with_reduction_147;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_148;
            end if;
        when square_with_reduction_148 => 
            next_state <= square_with_reduction_148;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_149;
            end if;
        when square_with_reduction_149 => 
            next_state <= square_with_reduction_149;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_150;
            end if;
        when square_with_reduction_150 => 
            next_state <= square_with_reduction_150;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_151;
            end if;
        when square_with_reduction_151 => 
            next_state <= square_with_reduction_151;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_152;
            end if;
        when square_with_reduction_152 => 
            next_state <= square_with_reduction_152;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_153;
            end if;
        when square_with_reduction_153 => 
            next_state <= square_with_reduction_153;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_154;
            end if;
        when square_with_reduction_154 => 
            next_state <= square_with_reduction_154;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_155;
            end if;
        when square_with_reduction_155 => 
            next_state <= square_with_reduction_155;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_156;
            end if;
        when square_with_reduction_156 => 
            next_state <= square_with_reduction_156;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_157;
            end if;
        when square_with_reduction_157 => 
            next_state <= square_with_reduction_157;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_158;
            end if;
        when square_with_reduction_158 => 
            next_state <= square_with_reduction_158;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_159;
            end if;
        when square_with_reduction_159 => 
            next_state <= square_with_reduction_159;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_160;
            end if;
        when square_with_reduction_160 => 
            next_state <= square_with_reduction_160;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_161;
            end if;
        when square_with_reduction_161 => 
            next_state <= square_with_reduction_161;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_162;
            end if;
        when square_with_reduction_162 => 
            next_state <= square_with_reduction_162;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_163;
            end if;
        when square_with_reduction_163 => 
            next_state <= square_with_reduction_163;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_164;
            end if;
        when square_with_reduction_164 => 
            next_state <= square_with_reduction_164;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_165;
            end if;
        when square_with_reduction_165 => 
            next_state <= square_with_reduction_165;
            if(penultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when square_with_reduction_167 => 
            next_state <= square_with_reduction_167;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_168;
            end if;
        when square_with_reduction_168 => 
            next_state <= square_with_reduction_168;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_169;
            end if;
        when square_with_reduction_169 => 
            next_state <= square_with_reduction_169;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_170;
            end if;
        when square_with_reduction_170 => 
            next_state <= square_with_reduction_170;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_171;
            end if;
        when square_with_reduction_171 => 
            next_state <= square_with_reduction_171;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_172;
            end if;
        when square_with_reduction_172 => 
            next_state <= square_with_reduction_172;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_173;
            end if;
        when square_with_reduction_173 => 
            next_state <= square_with_reduction_173;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_174;
            end if;
        when square_with_reduction_174 => 
            next_state <= square_with_reduction_174;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_175;
            end if;
        when square_with_reduction_175 => 
            next_state <= square_with_reduction_175;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_176;
            end if;
        when square_with_reduction_176 => 
            next_state <= square_with_reduction_176;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_177;
            end if;
        when square_with_reduction_177 => 
            next_state <= square_with_reduction_177;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_178;
            end if;
        when square_with_reduction_178 => 
            next_state <= square_with_reduction_178;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_179;
            end if;
        when square_with_reduction_179 => 
            next_state <= square_with_reduction_179;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_180;
            end if;
        when square_with_reduction_180 => 
            next_state <= square_with_reduction_180;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_181;
            end if;
        when square_with_reduction_181 => 
            next_state <= square_with_reduction_181;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_182;
            end if;
        when square_with_reduction_182 => 
            next_state <= square_with_reduction_182;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_183;
            end if;
        when square_with_reduction_183 => 
            next_state <= square_with_reduction_183;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_184;
            end if;
        when square_with_reduction_184 => 
            next_state <= square_with_reduction_184;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_185;
            end if;
        when square_with_reduction_185 => 
            next_state <= square_with_reduction_185;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_186;
            end if;
        when square_with_reduction_186 => 
            next_state <= square_with_reduction_186;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_187;
            end if;
        when square_with_reduction_187 => 
            next_state <= square_with_reduction_187;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_188;
            end if;
        when square_with_reduction_188 => 
            next_state <= square_with_reduction_188;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_189;
            end if;
        when square_with_reduction_189 => 
            next_state <= square_with_reduction_189;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_190;
            end if;
        when square_with_reduction_190 => 
            next_state <= square_with_reduction_190;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_191;
            end if;
        when square_with_reduction_191 => 
            next_state <= square_with_reduction_191;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_192;
            end if;
        when square_with_reduction_192 => 
            next_state <= square_with_reduction_192;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_193;
            end if;
        when square_with_reduction_193 => 
            next_state <= square_with_reduction_193;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_194;
            end if;
        when square_with_reduction_194 => 
            next_state <= square_with_reduction_194;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_195;
            end if;
        when square_with_reduction_195 => 
            next_state <= square_with_reduction_195;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_196;
            end if;
        when square_with_reduction_196 => 
            next_state <= square_with_reduction_196;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_197;
            end if;
        when square_with_reduction_197 => 
            next_state <= square_with_reduction_197;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_198;
            end if;
        when square_with_reduction_198 => 
            next_state <= square_with_reduction_198;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_199;
            end if;
        when square_with_reduction_199 => 
            next_state <= square_with_reduction_199;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_200;
            end if;
        when square_with_reduction_200 => 
            next_state <= square_with_reduction_200;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_201;
            end if;
        when square_with_reduction_201 => 
            next_state <= square_with_reduction_201;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_202;
            end if;
        when square_with_reduction_202 => 
            next_state <= square_with_reduction_202;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_203;
            end if;
        when square_with_reduction_203 => 
            next_state <= square_with_reduction_203;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_204;
            end if;
        when square_with_reduction_204 => 
            next_state <= square_with_reduction_204;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_205;
            end if;
        when square_with_reduction_205 => 
            next_state <= square_with_reduction_205;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_206;
            end if;
        when square_with_reduction_206 => 
            next_state <= square_with_reduction_206;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_207;
            end if;
        when square_with_reduction_207 => 
            next_state <= square_with_reduction_207;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_208;
            end if;
        when square_with_reduction_208 => 
            next_state <= square_with_reduction_208;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_209;
            end if;
        when square_with_reduction_209 => 
            next_state <= square_with_reduction_209;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_210;
            end if;
        when square_with_reduction_210 => 
            next_state <= square_with_reduction_210;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_211;
            end if;
        when square_with_reduction_211 => 
            next_state <= square_with_reduction_211;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_212;
            end if;
        when square_with_reduction_212 => 
            next_state <= square_with_reduction_212;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_213;
            end if;
        when square_with_reduction_213 => 
            next_state <= square_with_reduction_213;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_214;
            end if;
        when square_with_reduction_214 => 
            next_state <= square_with_reduction_214;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_215;
            end if;
        when square_with_reduction_215 => 
            next_state <= square_with_reduction_215;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_216;
            end if;
        when square_with_reduction_216 => 
            next_state <= square_with_reduction_216;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_217;
            end if;
        when square_with_reduction_217 => 
            next_state <= square_with_reduction_217;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_218;
            end if;
        when square_with_reduction_218 => 
            next_state <= square_with_reduction_218;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_219;
            end if;
        when square_with_reduction_219 => 
            next_state <= square_with_reduction_219;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_220;
            end if;
        when square_with_reduction_220 => 
            next_state <= square_with_reduction_220;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_221;
            end if;
        when square_with_reduction_221 => 
            next_state <= square_with_reduction_221;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_222;
            end if;
        when square_with_reduction_222 => 
            next_state <= square_with_reduction_222;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_223;
            end if;
        when square_with_reduction_223 => 
            next_state <= square_with_reduction_223;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_224;
            end if;
        when square_with_reduction_224 => 
            next_state <= square_with_reduction_224;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_225;
            end if;
        when square_with_reduction_225 => 
            next_state <= square_with_reduction_225;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_226;
            end if;
        when square_with_reduction_226 => 
            next_state <= square_with_reduction_226;
            if(penultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when square_with_reduction_special_prime_0 => 
            next_state <= square_with_reduction_special_prime_0;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1;
            end if;
        when square_with_reduction_special_prime_1 => 
            next_state <= square_with_reduction_special_prime_1;
            if(penultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when square_with_reduction_special_prime_3 => 
            next_state <= square_with_reduction_special_prime_3;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_4;
            end if;
        when square_with_reduction_special_prime_4 =>
            next_state <= square_with_reduction_special_prime_4;
            if(penultimate_operation = '1') then
                if(operands_size = "001") then
                    next_state <= square_with_reduction_special_prime_5;
                else
                    next_state <= square_with_reduction_special_prime_9;
                end if;
            end if;
        when square_with_reduction_special_prime_5 => 
            next_state <= square_with_reduction_special_prime_5;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_6;
            end if;
        when square_with_reduction_special_prime_6 => 
            next_state <= square_with_reduction_special_prime_6;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_7;
            end if;
        when square_with_reduction_special_prime_7 => 
            next_state <= square_with_reduction_special_prime_7;
            if(penultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when square_with_reduction_special_prime_9 => 
            next_state <= square_with_reduction_special_prime_9;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_10;
            end if;
        when square_with_reduction_special_prime_10 => 
            next_state <= square_with_reduction_special_prime_10;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_11;
            end if;
        when square_with_reduction_special_prime_11 => 
            next_state <= square_with_reduction_special_prime_11;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_12;
            end if;
        when square_with_reduction_special_prime_12 => 
            next_state <= square_with_reduction_special_prime_12;
            if(penultimate_operation = '1') then
                if(operands_size = "010") then
                    next_state <= square_with_reduction_special_prime_13;
                else
                    next_state <= square_with_reduction_special_prime_20;
                end if;
            end if;
        when square_with_reduction_special_prime_13 => 
            next_state <= square_with_reduction_special_prime_13;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_14;
            end if;
        when square_with_reduction_special_prime_14 => 
            next_state <= square_with_reduction_special_prime_14;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_15;
            end if;
        when square_with_reduction_special_prime_15 => 
            next_state <= square_with_reduction_special_prime_15;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_16;
            end if;
        when square_with_reduction_special_prime_16 => 
            next_state <= square_with_reduction_special_prime_16;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_17;
            end if;
        when square_with_reduction_special_prime_17 => 
            next_state <= square_with_reduction_special_prime_17;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_18;
            end if;
        when square_with_reduction_special_prime_18 => 
            next_state <= square_with_reduction_special_prime_18;
            if(penultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when square_with_reduction_special_prime_20 => 
            next_state <= square_with_reduction_special_prime_20;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_21;
            end if;
        when square_with_reduction_special_prime_21 => 
            next_state <= square_with_reduction_special_prime_21;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_22;
            end if;
        when square_with_reduction_special_prime_22 => 
            next_state <= square_with_reduction_special_prime_22;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_23;
            end if;
        when square_with_reduction_special_prime_23 => 
            next_state <= square_with_reduction_special_prime_23;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_24;
            end if;
        when square_with_reduction_special_prime_24 => 
            next_state <= square_with_reduction_special_prime_24;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_25;
            end if;
        when square_with_reduction_special_prime_25 => 
            next_state <= square_with_reduction_special_prime_25;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_26;
            end if;
        when square_with_reduction_special_prime_26 => 
            next_state <= square_with_reduction_special_prime_26;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_27;
            end if;
        when square_with_reduction_special_prime_27 => 
            next_state <= square_with_reduction_special_prime_27;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_28;
            end if;
        when square_with_reduction_special_prime_28 => 
            next_state <= square_with_reduction_special_prime_28;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_29;
            end if;
        when square_with_reduction_special_prime_29 => 
            next_state <= square_with_reduction_special_prime_29;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_30;
            end if;
        when square_with_reduction_special_prime_30 => 
            next_state <= square_with_reduction_special_prime_30;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_31;
            end if;
        when square_with_reduction_special_prime_31 => 
            next_state <= square_with_reduction_special_prime_31;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_32;
            end if;
        when square_with_reduction_special_prime_32 => 
            next_state <= square_with_reduction_special_prime_32;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_33;
            end if;
        when square_with_reduction_special_prime_33 => 
            next_state <= square_with_reduction_special_prime_33;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_34;
            end if;
        when square_with_reduction_special_prime_34 => 
            next_state <= square_with_reduction_special_prime_34;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_35;
            end if;
        when square_with_reduction_special_prime_35 => 
            next_state <= square_with_reduction_special_prime_35;
            if(penultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when square_with_reduction_special_prime_37 => 
            next_state <= square_with_reduction_special_prime_37;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_38;
            end if;
        when square_with_reduction_special_prime_38 => 
            next_state <= square_with_reduction_special_prime_38;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_39;
            end if;
        when square_with_reduction_special_prime_39 => 
            next_state <= square_with_reduction_special_prime_39;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_40;
            end if;
        when square_with_reduction_special_prime_40 => 
            next_state <= square_with_reduction_special_prime_40;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_41;
            end if;
        when square_with_reduction_special_prime_41 => 
            next_state <= square_with_reduction_special_prime_41;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_42;
            end if;
        when square_with_reduction_special_prime_42 => 
            next_state <= square_with_reduction_special_prime_42;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_43;
            end if;
        when square_with_reduction_special_prime_43 => 
            next_state <= square_with_reduction_special_prime_43;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_44;
            end if;
        when square_with_reduction_special_prime_44 => 
            next_state <= square_with_reduction_special_prime_44;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_45;
            end if;
        when square_with_reduction_special_prime_45 => 
            next_state <= square_with_reduction_special_prime_45;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_46;
            end if;
        when square_with_reduction_special_prime_46 => 
            next_state <= square_with_reduction_special_prime_46;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_47;
            end if;
        when square_with_reduction_special_prime_47 => 
            next_state <= square_with_reduction_special_prime_47;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_48;
            end if;
        when square_with_reduction_special_prime_48 => 
            next_state <= square_with_reduction_special_prime_48;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_49;
            end if;
        when square_with_reduction_special_prime_49 => 
            next_state <= square_with_reduction_special_prime_49;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_50;
            end if;
        when square_with_reduction_special_prime_50 => 
            next_state <= square_with_reduction_special_prime_50;
            if(penultimate_operation = '1') then
                if(operands_size = "100") then
                    next_state <= square_with_reduction_special_prime_51;
                else
                    next_state <= square_with_reduction_special_prime_68;
                end if;
            end if;
        when square_with_reduction_special_prime_51 => 
            next_state <= square_with_reduction_special_prime_51;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_52;
            end if;
        when square_with_reduction_special_prime_52 => 
            next_state <= square_with_reduction_special_prime_52;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_53;
            end if;
        when square_with_reduction_special_prime_53 => 
            next_state <= square_with_reduction_special_prime_53;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_54;
            end if;
        when square_with_reduction_special_prime_54 => 
            next_state <= square_with_reduction_special_prime_54;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_55;
            end if;
        when square_with_reduction_special_prime_55 => 
            next_state <= square_with_reduction_special_prime_55;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_56;
            end if;
        when square_with_reduction_special_prime_56 => 
            next_state <= square_with_reduction_special_prime_56;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_57;
            end if;
        when square_with_reduction_special_prime_57 => 
            next_state <= square_with_reduction_special_prime_57;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_58;
            end if;
        when square_with_reduction_special_prime_58 => 
            next_state <= square_with_reduction_special_prime_58;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_59;
            end if;
        when square_with_reduction_special_prime_59 => 
            next_state <= square_with_reduction_special_prime_59;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_60;
            end if;
        when square_with_reduction_special_prime_60 => 
            next_state <= square_with_reduction_special_prime_60;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_61;
            end if;
        when square_with_reduction_special_prime_61 => 
            next_state <= square_with_reduction_special_prime_61;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_62;
            end if;
        when square_with_reduction_special_prime_62 => 
            next_state <= square_with_reduction_special_prime_62;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_63;
            end if;
        when square_with_reduction_special_prime_63 => 
            next_state <= square_with_reduction_special_prime_63;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_64;
            end if;
        when square_with_reduction_special_prime_64 => 
            next_state <= square_with_reduction_special_prime_64;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_65;
            end if;
        when square_with_reduction_special_prime_65 => 
            next_state <= square_with_reduction_special_prime_65;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_66;
            end if;
        when square_with_reduction_special_prime_66 => 
            next_state <= square_with_reduction_special_prime_66;
            if(penultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when square_with_reduction_special_prime_68 => 
            next_state <= square_with_reduction_special_prime_68;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_69;
            end if;
        when square_with_reduction_special_prime_69 => 
            next_state <= square_with_reduction_special_prime_69;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_70;
            end if;
        when square_with_reduction_special_prime_70 => 
            next_state <= square_with_reduction_special_prime_70;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_71;
            end if;
        when square_with_reduction_special_prime_71 => 
            next_state <= square_with_reduction_special_prime_71;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_72;
            end if;
        when square_with_reduction_special_prime_72 => 
            next_state <= square_with_reduction_special_prime_72;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_73;
            end if;
        when square_with_reduction_special_prime_73 => 
            next_state <= square_with_reduction_special_prime_73;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_74;
            end if;
        when square_with_reduction_special_prime_74 => 
            next_state <= square_with_reduction_special_prime_74;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_75;
            end if;
        when square_with_reduction_special_prime_75 => 
            next_state <= square_with_reduction_special_prime_75;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_76;
            end if;
        when square_with_reduction_special_prime_76 => 
            next_state <= square_with_reduction_special_prime_76;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_77;
            end if;
        when square_with_reduction_special_prime_77 => 
            next_state <= square_with_reduction_special_prime_77;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_78;
            end if;
        when square_with_reduction_special_prime_78 => 
            next_state <= square_with_reduction_special_prime_78;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_79;
            end if;
        when square_with_reduction_special_prime_79 => 
            next_state <= square_with_reduction_special_prime_79;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_80;
            end if;
        when square_with_reduction_special_prime_80 => 
            next_state <= square_with_reduction_special_prime_80;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_81;
            end if;
        when square_with_reduction_special_prime_81 => 
            next_state <= square_with_reduction_special_prime_81;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_82;
            end if;
        when square_with_reduction_special_prime_82 => 
            next_state <= square_with_reduction_special_prime_82;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_83;
            end if;
        when square_with_reduction_special_prime_83 => 
            next_state <= square_with_reduction_special_prime_83;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_84;
            end if;
        when square_with_reduction_special_prime_84 => 
            next_state <= square_with_reduction_special_prime_84;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_85;
            end if;
        when square_with_reduction_special_prime_85 => 
            next_state <= square_with_reduction_special_prime_85;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_86;
            end if;
        when square_with_reduction_special_prime_86 => 
            next_state <= square_with_reduction_special_prime_86;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_87;
            end if;
        when square_with_reduction_special_prime_87 => 
            next_state <= square_with_reduction_special_prime_87;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_88;
            end if;
        when square_with_reduction_special_prime_88 => 
            next_state <= square_with_reduction_special_prime_88;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_89;
            end if;
        when square_with_reduction_special_prime_89 => 
            next_state <= square_with_reduction_special_prime_89;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_90;
            end if;
        when square_with_reduction_special_prime_90 => 
            next_state <= square_with_reduction_special_prime_90;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_91;
            end if;
        when square_with_reduction_special_prime_91 => 
            next_state <= square_with_reduction_special_prime_91;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_92;
            end if;
        when square_with_reduction_special_prime_92 => 
            next_state <= square_with_reduction_special_prime_92;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_93;
            end if;
        when square_with_reduction_special_prime_93 => 
            next_state <= square_with_reduction_special_prime_93;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_94;
            end if;
        when square_with_reduction_special_prime_94 => 
            next_state <= square_with_reduction_special_prime_94;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_95;
            end if;
        when square_with_reduction_special_prime_95 => 
            next_state <= square_with_reduction_special_prime_95;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_96;
            end if;
        when square_with_reduction_special_prime_96 => 
            next_state <= square_with_reduction_special_prime_96;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_97;
            end if;
        when square_with_reduction_special_prime_97 => 
            next_state <= square_with_reduction_special_prime_97;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_98;
            end if;
        when square_with_reduction_special_prime_98 => 
            next_state <= square_with_reduction_special_prime_98;
            if(penultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when square_with_reduction_special_prime_100 => 
            next_state <= square_with_reduction_special_prime_100;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_101;
            end if;
        when square_with_reduction_special_prime_101 => 
            next_state <= square_with_reduction_special_prime_101;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_102;
            end if;
        when square_with_reduction_special_prime_102 => 
            next_state <= square_with_reduction_special_prime_102;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_103;
            end if;
        when square_with_reduction_special_prime_103 => 
            next_state <= square_with_reduction_special_prime_103;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_104;
            end if;
        when square_with_reduction_special_prime_104 => 
            next_state <= square_with_reduction_special_prime_104;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_105;
            end if;
        when square_with_reduction_special_prime_105 => 
            next_state <= square_with_reduction_special_prime_105;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_106;
            end if;
        when square_with_reduction_special_prime_106 => 
            next_state <= square_with_reduction_special_prime_106;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_107;
            end if;
        when square_with_reduction_special_prime_107 => 
            next_state <= square_with_reduction_special_prime_107;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_108;
            end if;
        when square_with_reduction_special_prime_108 => 
            next_state <= square_with_reduction_special_prime_108;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_109;
            end if;
        when square_with_reduction_special_prime_109 => 
            next_state <= square_with_reduction_special_prime_109;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_110;
            end if;
        when square_with_reduction_special_prime_110 => 
            next_state <= square_with_reduction_special_prime_110;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_111;
            end if;
        when square_with_reduction_special_prime_111 => 
            next_state <= square_with_reduction_special_prime_111;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_112;
            end if;
        when square_with_reduction_special_prime_112 => 
            next_state <= square_with_reduction_special_prime_112;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_113;
            end if;
        when square_with_reduction_special_prime_113 => 
            next_state <= square_with_reduction_special_prime_113;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_114;
            end if;
        when square_with_reduction_special_prime_114 => 
            next_state <= square_with_reduction_special_prime_114;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_115;
            end if;
        when square_with_reduction_special_prime_115 => 
            next_state <= square_with_reduction_special_prime_115;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_116;
            end if;
        when square_with_reduction_special_prime_116 => 
            next_state <= square_with_reduction_special_prime_116;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_117;
            end if;
        when square_with_reduction_special_prime_117 => 
            next_state <= square_with_reduction_special_prime_117;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_118;
            end if;
        when square_with_reduction_special_prime_118 => 
            next_state <= square_with_reduction_special_prime_118;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_119;
            end if;
        when square_with_reduction_special_prime_119 => 
            next_state <= square_with_reduction_special_prime_119;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_120;
            end if;
        when square_with_reduction_special_prime_120 => 
            next_state <= square_with_reduction_special_prime_120;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_121;
            end if;
        when square_with_reduction_special_prime_121 => 
            next_state <= square_with_reduction_special_prime_121;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_122;
            end if;
        when square_with_reduction_special_prime_122 => 
            next_state <= square_with_reduction_special_prime_122;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_123;
            end if;
        when square_with_reduction_special_prime_123 => 
            next_state <= square_with_reduction_special_prime_123;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_124;
            end if;
        when square_with_reduction_special_prime_124 => 
            next_state <= square_with_reduction_special_prime_124;
            if(penultimate_operation = '1') then
                if(operands_size = "110") then
                    next_state <= square_with_reduction_special_prime_125;
                else
                    next_state <= square_with_reduction_special_prime_157;
                end if;
            end if;
        when square_with_reduction_special_prime_125 => 
            next_state <= square_with_reduction_special_prime_125;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_126;
            end if;
        when square_with_reduction_special_prime_126 => 
            next_state <= square_with_reduction_special_prime_126;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_127;
            end if;
        when square_with_reduction_special_prime_127 => 
            next_state <= square_with_reduction_special_prime_127;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_128;
            end if;
        when square_with_reduction_special_prime_128 => 
            next_state <= square_with_reduction_special_prime_128;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_129;
            end if;
        when square_with_reduction_special_prime_129 => 
            next_state <= square_with_reduction_special_prime_129;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_130;
            end if;
        when square_with_reduction_special_prime_130 => 
            next_state <= square_with_reduction_special_prime_130;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_131;
            end if;
        when square_with_reduction_special_prime_131 => 
            next_state <= square_with_reduction_special_prime_131;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_132;
            end if;
        when square_with_reduction_special_prime_132 => 
            next_state <= square_with_reduction_special_prime_132;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_133;
            end if;
        when square_with_reduction_special_prime_133 => 
            next_state <= square_with_reduction_special_prime_133;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_134;
            end if;
        when square_with_reduction_special_prime_134 => 
            next_state <= square_with_reduction_special_prime_134;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_135;
            end if;
        when square_with_reduction_special_prime_135 => 
            next_state <= square_with_reduction_special_prime_135;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_136;
            end if;
        when square_with_reduction_special_prime_136 => 
            next_state <= square_with_reduction_special_prime_136;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_137;
            end if;
        when square_with_reduction_special_prime_137 => 
            next_state <= square_with_reduction_special_prime_137;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_138;
            end if;
        when square_with_reduction_special_prime_138 => 
            next_state <= square_with_reduction_special_prime_138;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_139;
            end if;
        when square_with_reduction_special_prime_139 => 
            next_state <= square_with_reduction_special_prime_139;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_140;
            end if;
        when square_with_reduction_special_prime_140 => 
            next_state <= square_with_reduction_special_prime_140;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_141;
            end if;
        when square_with_reduction_special_prime_141 => 
            next_state <= square_with_reduction_special_prime_141;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_142;
            end if;
        when square_with_reduction_special_prime_142 => 
            next_state <= square_with_reduction_special_prime_142;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_143;
            end if;
        when square_with_reduction_special_prime_143 => 
            next_state <= square_with_reduction_special_prime_143;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_144;
            end if;
        when square_with_reduction_special_prime_144 => 
            next_state <= square_with_reduction_special_prime_144;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_145;
            end if;
        when square_with_reduction_special_prime_145 => 
            next_state <= square_with_reduction_special_prime_145;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_146;
            end if;
        when square_with_reduction_special_prime_146 => 
            next_state <= square_with_reduction_special_prime_146;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_147;
            end if;
        when square_with_reduction_special_prime_147 => 
            next_state <= square_with_reduction_special_prime_147;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_148;
            end if;
        when square_with_reduction_special_prime_148 => 
            next_state <= square_with_reduction_special_prime_148;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_149;
            end if;
        when square_with_reduction_special_prime_149 => 
            next_state <= square_with_reduction_special_prime_149;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_150;
            end if;
        when square_with_reduction_special_prime_150 => 
            next_state <= square_with_reduction_special_prime_150;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_151;
            end if;
        when square_with_reduction_special_prime_151 => 
            next_state <= square_with_reduction_special_prime_151;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_152;
            end if;
        when square_with_reduction_special_prime_152 => 
            next_state <= square_with_reduction_special_prime_152;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_153;
            end if;
        when square_with_reduction_special_prime_153 => 
            next_state <= square_with_reduction_special_prime_153;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_154;
            end if;
        when square_with_reduction_special_prime_154 => 
            next_state <= square_with_reduction_special_prime_154;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_155;
            end if;            
        when square_with_reduction_special_prime_155 => 
            next_state <= square_with_reduction_special_prime_155;
            if(penultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when square_with_reduction_special_prime_157 => 
            next_state <= square_with_reduction_special_prime_157;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_158;
            end if;
        when square_with_reduction_special_prime_158 => 
            next_state <= square_with_reduction_special_prime_158;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_159;
            end if;
        when square_with_reduction_special_prime_159 => 
            next_state <= square_with_reduction_special_prime_159;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_160;
            end if;
        when square_with_reduction_special_prime_160 => 
            next_state <= square_with_reduction_special_prime_160;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_161;
            end if;
        when square_with_reduction_special_prime_161 => 
            next_state <= square_with_reduction_special_prime_161;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_162;
            end if;
        when square_with_reduction_special_prime_162 => 
            next_state <= square_with_reduction_special_prime_162;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_163;
            end if;
        when square_with_reduction_special_prime_163 => 
            next_state <= square_with_reduction_special_prime_163;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_164;
            end if;
        when square_with_reduction_special_prime_164 => 
            next_state <= square_with_reduction_special_prime_164;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_165;
            end if;
        when square_with_reduction_special_prime_165 => 
            next_state <= square_with_reduction_special_prime_165;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_166;
            end if;
        when square_with_reduction_special_prime_166 => 
            next_state <= square_with_reduction_special_prime_166;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_167;
            end if;
        when square_with_reduction_special_prime_167 => 
            next_state <= square_with_reduction_special_prime_167;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_168;
            end if;
        when square_with_reduction_special_prime_168 => 
            next_state <= square_with_reduction_special_prime_168;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_169;
            end if;
        when square_with_reduction_special_prime_169 => 
            next_state <= square_with_reduction_special_prime_169;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_170;
            end if;
        when square_with_reduction_special_prime_170 => 
            next_state <= square_with_reduction_special_prime_170;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_171;
            end if;
        when square_with_reduction_special_prime_171 => 
            next_state <= square_with_reduction_special_prime_171;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_172;
            end if;
        when square_with_reduction_special_prime_172 => 
            next_state <= square_with_reduction_special_prime_172;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_173;
            end if;
        when square_with_reduction_special_prime_173 => 
            next_state <= square_with_reduction_special_prime_173;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_174;
            end if;
        when square_with_reduction_special_prime_174 => 
            next_state <= square_with_reduction_special_prime_174;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_175;
            end if;
        when square_with_reduction_special_prime_175 => 
            next_state <= square_with_reduction_special_prime_175;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_176;
            end if;
        when square_with_reduction_special_prime_176 => 
            next_state <= square_with_reduction_special_prime_176;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_177;
            end if;
        when square_with_reduction_special_prime_177 => 
            next_state <= square_with_reduction_special_prime_177;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_178;
            end if;
        when square_with_reduction_special_prime_178 => 
            next_state <= square_with_reduction_special_prime_178;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_179;
            end if;
        when square_with_reduction_special_prime_179 => 
            next_state <= square_with_reduction_special_prime_179;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_180;
            end if;
        when square_with_reduction_special_prime_180 => 
            next_state <= square_with_reduction_special_prime_180;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_181;
            end if;
        when square_with_reduction_special_prime_181 => 
            next_state <= square_with_reduction_special_prime_181;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_182;
            end if;
        when square_with_reduction_special_prime_182 => 
            next_state <= square_with_reduction_special_prime_182;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_183;
            end if;
        when square_with_reduction_special_prime_183 => 
            next_state <= square_with_reduction_special_prime_183;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_184;
            end if;
        when square_with_reduction_special_prime_184 => 
            next_state <= square_with_reduction_special_prime_184;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_185;
            end if;
        when square_with_reduction_special_prime_185 => 
            next_state <= square_with_reduction_special_prime_185;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_186;
            end if;
        when square_with_reduction_special_prime_186 => 
            next_state <= square_with_reduction_special_prime_186;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_187;
            end if;
        when square_with_reduction_special_prime_187 => 
            next_state <= square_with_reduction_special_prime_187;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_188;
            end if;
        when square_with_reduction_special_prime_188 => 
            next_state <= square_with_reduction_special_prime_188;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_189;
            end if;
        when square_with_reduction_special_prime_189 => 
            next_state <= square_with_reduction_special_prime_189;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_190;
            end if;
        when square_with_reduction_special_prime_190 => 
            next_state <= square_with_reduction_special_prime_190;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_191;
            end if;
        when square_with_reduction_special_prime_191 => 
            next_state <= square_with_reduction_special_prime_191;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_192;
            end if;
        when square_with_reduction_special_prime_192 => 
            next_state <= square_with_reduction_special_prime_192;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_193;
            end if;
        when square_with_reduction_special_prime_193 => 
            next_state <= square_with_reduction_special_prime_193;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_194;
            end if;
        when square_with_reduction_special_prime_194 => 
            next_state <= square_with_reduction_special_prime_194;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_195;
            end if;
        when square_with_reduction_special_prime_195 => 
            next_state <= square_with_reduction_special_prime_195;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_196;
            end if;
        when square_with_reduction_special_prime_196 => 
            next_state <= square_with_reduction_special_prime_196;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_197;
            end if;
        when square_with_reduction_special_prime_197 => 
            next_state <= square_with_reduction_special_prime_197;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_198;
            end if;
        when square_with_reduction_special_prime_198 => 
            next_state <= square_with_reduction_special_prime_198;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_199;
            end if;
        when square_with_reduction_special_prime_199 => 
            next_state <= square_with_reduction_special_prime_199;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_200;
            end if;
        when square_with_reduction_special_prime_200 => 
            next_state <= square_with_reduction_special_prime_200;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_201;
            end if;
        when square_with_reduction_special_prime_201 => 
            next_state <= square_with_reduction_special_prime_201;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_202;
            end if;
        when square_with_reduction_special_prime_202 => 
            next_state <= square_with_reduction_special_prime_202;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_203;
            end if;
        when square_with_reduction_special_prime_203 => 
            next_state <= square_with_reduction_special_prime_203;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_204;
            end if;
        when square_with_reduction_special_prime_204 => 
            next_state <= square_with_reduction_special_prime_204;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_205;
            end if;
        when square_with_reduction_special_prime_205 => 
            next_state <= square_with_reduction_special_prime_205;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_206;
            end if;
        when square_with_reduction_special_prime_206 => 
            next_state <= square_with_reduction_special_prime_206;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_207;
            end if;
        when square_with_reduction_special_prime_207 => 
            next_state <= square_with_reduction_special_prime_207;
            if(penultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when addition_subtraction_direct_0 =>
            next_state <= addition_subtraction_direct_0;
            if(penultimate_operation = '1') then
                next_state <= nop_4_stages;
            end if;
        when addition_subtraction_direct_2 =>
            next_state <= addition_subtraction_direct_2;
            if(penultimate_operation = '1') then
                if(operands_size = "001") then
                    next_state <= addition_subtraction_direct_3;
                else
                    next_state <= addition_subtraction_direct_5;
                end if;
            end if;
        when addition_subtraction_direct_3 =>
            next_state <= addition_subtraction_direct_3;
            if(penultimate_operation = '1') then
                next_state <= nop_4_stages;
            end if;
        when addition_subtraction_direct_5 =>
            next_state <= addition_subtraction_direct_5;
            if(penultimate_operation = '1') then
                if(operands_size = "010") then
                    next_state <= addition_subtraction_direct_6;
                else
                    next_state <= addition_subtraction_direct_8;
                end if;
            end if;
        when addition_subtraction_direct_6 =>
            next_state <= addition_subtraction_direct_6;
            if(penultimate_operation = '1') then
                next_state <= nop_4_stages;
            end if;
        when addition_subtraction_direct_8 =>
            next_state <= addition_subtraction_direct_8;
            if(penultimate_operation = '1') then
                if(operands_size = "011") then
                    next_state <= addition_subtraction_direct_9;
                else
                    next_state <= addition_subtraction_direct_11;
                end if;
            end if;
        when addition_subtraction_direct_9 =>
            next_state <= addition_subtraction_direct_9;
            if(penultimate_operation = '1') then
                next_state <= nop_4_stages;
            end if;
        when addition_subtraction_direct_11 =>
            next_state <= addition_subtraction_direct_11;
            if(penultimate_operation = '1') then
                if(operands_size = "100") then
                    next_state <= addition_subtraction_direct_12;
                else
                    next_state <= addition_subtraction_direct_14;
                end if;
            end if;
        when addition_subtraction_direct_12 =>
            next_state <= addition_subtraction_direct_12;
            if(penultimate_operation = '1') then
                next_state <= nop_4_stages;
            end if;
        when addition_subtraction_direct_14 =>
            next_state <= addition_subtraction_direct_14;
            if(penultimate_operation = '1') then
                if(operands_size = "101") then
                    next_state <= addition_subtraction_direct_15;
                else
                    next_state <= addition_subtraction_direct_17;
                end if;
            end if;
        when addition_subtraction_direct_15 =>
            next_state <= addition_subtraction_direct_15;
            if(penultimate_operation = '1') then
                next_state <= nop_4_stages;
            end if;
        when addition_subtraction_direct_17 =>
            next_state <= addition_subtraction_direct_17;
            if(penultimate_operation = '1') then
                if(operands_size = "110") then
                    next_state <= addition_subtraction_direct_18;
                else
                    next_state <= addition_subtraction_direct_20;
                end if;
            end if;
        when addition_subtraction_direct_18 =>
            next_state <= addition_subtraction_direct_18;
            if(penultimate_operation = '1') then
                next_state <= nop_4_stages;
            end if;
        when addition_subtraction_direct_20 =>
            next_state <= addition_subtraction_direct_20;
            if(penultimate_operation = '1') then
                next_state <= addition_subtraction_direct_21;
            end if;
        when addition_subtraction_direct_21 =>
            next_state <= addition_subtraction_direct_21;
            if(penultimate_operation = '1') then
                next_state <= nop_4_stages;
            end if;
        when iterative_modular_reduction_0 =>
            next_state <= iterative_modular_reduction_0;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_1;
            end if;    
        when iterative_modular_reduction_1 =>
            next_state <= iterative_modular_reduction_1;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_2;
            end if;
        when iterative_modular_reduction_2 =>
            next_state <= iterative_modular_reduction_2;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_3;
            end if;
        when iterative_modular_reduction_3 =>
            next_state <= iterative_modular_reduction_3;
            if(penultimate_operation = '1') then
                next_state <= nop_4_stages;
            end if;
        when iterative_modular_reduction_5 =>
            next_state <= iterative_modular_reduction_5;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_6;
            end if;
        when iterative_modular_reduction_6 =>
            next_state <= iterative_modular_reduction_6;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_7;
            end if;
        when iterative_modular_reduction_7 =>
            next_state <= iterative_modular_reduction_7;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_8;
            end if;
        when iterative_modular_reduction_8 =>
            next_state <= iterative_modular_reduction_8;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_9;
            end if;
        when iterative_modular_reduction_9 =>
            next_state <= iterative_modular_reduction_9;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_10;
            end if;
        when iterative_modular_reduction_10 =>
            next_state <= iterative_modular_reduction_10;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_11;
            end if;
        when iterative_modular_reduction_11 =>
            next_state <= iterative_modular_reduction_11;
            if(penultimate_operation = '1') then
                next_state <= nop_4_stages;
            end if;
        when iterative_modular_reduction_13 =>
            next_state <= iterative_modular_reduction_13;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_14;
            end if;
        when iterative_modular_reduction_14 =>
            next_state <= iterative_modular_reduction_14;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_15;
            end if;
        when iterative_modular_reduction_15 =>
            next_state <= iterative_modular_reduction_15;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_16;
            end if;
        when iterative_modular_reduction_16 =>
            next_state <= iterative_modular_reduction_16;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_17;
            end if;
        when iterative_modular_reduction_17 =>
            next_state <= iterative_modular_reduction_17;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_18;
            end if;
        when iterative_modular_reduction_18 =>
            next_state <= iterative_modular_reduction_18;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_19;
            end if;
        when iterative_modular_reduction_19 =>
            next_state <= iterative_modular_reduction_19;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_20;
            end if;
        when iterative_modular_reduction_20 =>
            next_state <= iterative_modular_reduction_20;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_21;
            end if;
        when iterative_modular_reduction_21 =>
            next_state <= iterative_modular_reduction_21;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_22;
            end if;
        when iterative_modular_reduction_22 =>
            next_state <= iterative_modular_reduction_22;
            if(penultimate_operation = '1') then
                next_state <= nop_4_stages;
            end if;
        when iterative_modular_reduction_24 =>
            next_state <= iterative_modular_reduction_24;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_25;
            end if;
        when iterative_modular_reduction_25 =>
            next_state <= iterative_modular_reduction_25;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_26;
            end if;
        when iterative_modular_reduction_26 =>
            next_state <= iterative_modular_reduction_26;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_27;
            end if;
        when iterative_modular_reduction_27 =>
            next_state <= iterative_modular_reduction_27;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_28;
            end if;
        when iterative_modular_reduction_28 =>
            next_state <= iterative_modular_reduction_28;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_29;
            end if;
        when iterative_modular_reduction_29 =>
            next_state <= iterative_modular_reduction_29;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_30;
            end if;
        when iterative_modular_reduction_30 =>
            next_state <= iterative_modular_reduction_30;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_31;
            end if;
        when iterative_modular_reduction_31 =>
            next_state <= iterative_modular_reduction_31;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_32;
            end if;
        when iterative_modular_reduction_32 =>
            next_state <= iterative_modular_reduction_32;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_33;
            end if;
        when iterative_modular_reduction_33 =>
            next_state <= iterative_modular_reduction_33;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_34;
            end if;
        when iterative_modular_reduction_34 =>
            next_state <= iterative_modular_reduction_34;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_35;
            end if;
        when iterative_modular_reduction_35 =>
            next_state <= iterative_modular_reduction_35;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_36;
            end if;
        when iterative_modular_reduction_36 =>
            next_state <= iterative_modular_reduction_36;
            if(penultimate_operation = '1') then
                next_state <= nop_4_stages;
            end if;
        when iterative_modular_reduction_38 =>
            next_state <= iterative_modular_reduction_38;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_39;
            end if;
        when iterative_modular_reduction_39 =>
            next_state <= iterative_modular_reduction_39;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_40;
            end if;
        when iterative_modular_reduction_40 =>
            next_state <= iterative_modular_reduction_40;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_41;
            end if;
        when iterative_modular_reduction_41 =>
            next_state <= iterative_modular_reduction_41;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_42;
            end if;
        when iterative_modular_reduction_42 =>
            next_state <= iterative_modular_reduction_42;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_43;
            end if;
        when iterative_modular_reduction_43 =>
            next_state <= iterative_modular_reduction_43;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_44;
            end if;
        when iterative_modular_reduction_44 =>
            next_state <= iterative_modular_reduction_44;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_45;
            end if;
        when iterative_modular_reduction_45 =>
            next_state <= iterative_modular_reduction_45;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_46;
            end if;
        when iterative_modular_reduction_46 =>
            next_state <= iterative_modular_reduction_46;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_47;
            end if;
        when iterative_modular_reduction_47 =>
            next_state <= iterative_modular_reduction_47;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_48;
            end if;
        when iterative_modular_reduction_48 =>
            next_state <= iterative_modular_reduction_48;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_49;
            end if;
        when iterative_modular_reduction_49 =>
            next_state <= iterative_modular_reduction_49;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_50;
            end if;
        when iterative_modular_reduction_50 =>
            next_state <= iterative_modular_reduction_50;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_51;
            end if;
        when iterative_modular_reduction_51 =>
            next_state <= iterative_modular_reduction_51;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_52;
            end if;
        when iterative_modular_reduction_52 =>
            next_state <= iterative_modular_reduction_52;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_53;
            end if;
        when iterative_modular_reduction_53 =>
            next_state <= iterative_modular_reduction_53;
            if(penultimate_operation = '1') then
                next_state <= nop_4_stages;
            end if;
        when iterative_modular_reduction_55 =>
            next_state <= iterative_modular_reduction_55;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_56;
            end if;
        when iterative_modular_reduction_56 =>
            next_state <= iterative_modular_reduction_56;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_57;
            end if;
        when iterative_modular_reduction_57 =>
            next_state <= iterative_modular_reduction_57;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_58;
            end if;
        when iterative_modular_reduction_58 =>
            next_state <= iterative_modular_reduction_58;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_59;
            end if;
        when iterative_modular_reduction_59 =>
            next_state <= iterative_modular_reduction_59;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_60;
            end if;
        when iterative_modular_reduction_60 =>
            next_state <= iterative_modular_reduction_60;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_61;
            end if;
        when iterative_modular_reduction_61 =>
            next_state <= iterative_modular_reduction_61;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_62;
            end if;
        when iterative_modular_reduction_62 =>
            next_state <= iterative_modular_reduction_62;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_63;
            end if;
        when iterative_modular_reduction_63 =>
            next_state <= iterative_modular_reduction_63;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_64;
            end if;
        when iterative_modular_reduction_64 =>
            next_state <= iterative_modular_reduction_64;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_65;
            end if;
        when iterative_modular_reduction_65 =>
            next_state <= iterative_modular_reduction_65;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_66;
            end if;
        when iterative_modular_reduction_66 =>
            next_state <= iterative_modular_reduction_66;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_67;
            end if;
        when iterative_modular_reduction_67 =>
            next_state <= iterative_modular_reduction_67;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_68;
            end if;
        when iterative_modular_reduction_68 =>
            next_state <= iterative_modular_reduction_68;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_69;
            end if;
        when iterative_modular_reduction_69 =>
            next_state <= iterative_modular_reduction_69;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_70;
            end if;
        when iterative_modular_reduction_70 =>
            next_state <= iterative_modular_reduction_70;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_71;
            end if;
        when iterative_modular_reduction_71 =>
            next_state <= iterative_modular_reduction_71;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_72;
            end if;
        when iterative_modular_reduction_72 =>
            next_state <= iterative_modular_reduction_72;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_73;
            end if;
        when iterative_modular_reduction_73 =>
            next_state <= iterative_modular_reduction_73;
            if(penultimate_operation = '1') then
                next_state <= nop_4_stages;
            end if;
        when iterative_modular_reduction_75 =>
            next_state <= iterative_modular_reduction_75;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_76;
            end if;
        when iterative_modular_reduction_76 =>
            next_state <= iterative_modular_reduction_76;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_77;
            end if;
        when iterative_modular_reduction_77 =>
            next_state <= iterative_modular_reduction_77;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_78;
            end if;
        when iterative_modular_reduction_78 =>
            next_state <= iterative_modular_reduction_78;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_79;
            end if;
        when iterative_modular_reduction_79 =>
            next_state <= iterative_modular_reduction_79;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_80;
            end if;
        when iterative_modular_reduction_80 =>
            next_state <= iterative_modular_reduction_80;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_81;
            end if;
        when iterative_modular_reduction_81 =>
            next_state <= iterative_modular_reduction_81;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_82;
            end if;
        when iterative_modular_reduction_82 =>
            next_state <= iterative_modular_reduction_82;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_83;
            end if;
        when iterative_modular_reduction_83 =>
            next_state <= iterative_modular_reduction_83;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_84;
            end if;
        when iterative_modular_reduction_84 =>
            next_state <= iterative_modular_reduction_84;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_85;
            end if;
        when iterative_modular_reduction_85 =>
            next_state <= iterative_modular_reduction_85;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_86;
            end if;
        when iterative_modular_reduction_86 =>
            next_state <= iterative_modular_reduction_86;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_87;
            end if;
        when iterative_modular_reduction_87 =>
            next_state <= iterative_modular_reduction_87;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_88;
            end if;
        when iterative_modular_reduction_88 =>
            next_state <= iterative_modular_reduction_88;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_89;
            end if;
        when iterative_modular_reduction_89 =>
            next_state <= iterative_modular_reduction_89;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_90;
            end if;
        when iterative_modular_reduction_90 =>
            next_state <= iterative_modular_reduction_90;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_91;
            end if;
        when iterative_modular_reduction_91 =>
            next_state <= iterative_modular_reduction_91;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_92;
            end if;
        when iterative_modular_reduction_92 =>
            next_state <= iterative_modular_reduction_92;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_93;
            end if;
        when iterative_modular_reduction_93 =>
            next_state <= iterative_modular_reduction_93;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_94;
            end if;
        when iterative_modular_reduction_94 =>
            next_state <= iterative_modular_reduction_94;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_95;
            end if;
        when iterative_modular_reduction_95 =>
            next_state <= iterative_modular_reduction_95;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_96;
            end if;
        when iterative_modular_reduction_96 =>
            next_state <= iterative_modular_reduction_96;
            if(penultimate_operation = '1') then
                next_state <= nop_4_stages;
            end if;
        when iterative_modular_reduction_98 =>
            next_state <= iterative_modular_reduction_98;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_99;
            end if;
        when iterative_modular_reduction_99 =>
            next_state <= iterative_modular_reduction_99;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_100;
            end if;
        when iterative_modular_reduction_100 =>
            next_state <= iterative_modular_reduction_100;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_101;
            end if;
        when iterative_modular_reduction_101 =>
            next_state <= iterative_modular_reduction_101;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_102;
            end if;
        when iterative_modular_reduction_102 =>
            next_state <= iterative_modular_reduction_102;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_103;
            end if;
        when iterative_modular_reduction_103 =>
            next_state <= iterative_modular_reduction_103;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_104;
            end if;
        when iterative_modular_reduction_104 =>
            next_state <= iterative_modular_reduction_104;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_105;
            end if;
        when iterative_modular_reduction_105 =>
            next_state <= iterative_modular_reduction_105;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_106;
            end if;
        when iterative_modular_reduction_106 =>
            next_state <= iterative_modular_reduction_106;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_107;
            end if;
        when iterative_modular_reduction_107 =>
            next_state <= iterative_modular_reduction_107;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_108;
            end if;
        when iterative_modular_reduction_108 =>
            next_state <= iterative_modular_reduction_108;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_109;
            end if;
        when iterative_modular_reduction_109 =>
            next_state <= iterative_modular_reduction_109;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_110;
            end if;
        when iterative_modular_reduction_110 =>
            next_state <= iterative_modular_reduction_110;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_111;
            end if;
        when iterative_modular_reduction_111 =>
            next_state <= iterative_modular_reduction_111;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_112;
            end if;
        when iterative_modular_reduction_112 =>
            next_state <= iterative_modular_reduction_112;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_113;
            end if;
        when iterative_modular_reduction_113 =>
            next_state <= iterative_modular_reduction_113;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_114;
            end if;
        when iterative_modular_reduction_114 =>
            next_state <= iterative_modular_reduction_114;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_115;
            end if;
        when iterative_modular_reduction_115 =>
            next_state <= iterative_modular_reduction_115;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_116;
            end if;
        when iterative_modular_reduction_116 =>
            next_state <= iterative_modular_reduction_116;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_117;
            end if;
        when iterative_modular_reduction_117 =>
            next_state <= iterative_modular_reduction_117;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_118;
            end if;
        when iterative_modular_reduction_118 =>
            next_state <= iterative_modular_reduction_118;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_119;
            end if;
        when iterative_modular_reduction_119 =>
            next_state <= iterative_modular_reduction_119;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_120;
            end if;
        when iterative_modular_reduction_120 =>
            next_state <= iterative_modular_reduction_120;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_121;
            end if;
        when iterative_modular_reduction_121 =>
            next_state <= iterative_modular_reduction_121;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_122;
            end if;
        when iterative_modular_reduction_122 =>
            next_state <= iterative_modular_reduction_122;
            if(penultimate_operation = '1') then
                next_state <= nop_4_stages;
            end if;
        when nop_4_stages =>
            next_state <= nop_4_stages;
            if(penultimate_operation = '1') then
                next_state <= decode_instruction;
            end if;
        when nop_8_stages =>
            next_state <= nop_8_stages;
            if(penultimate_operation = '1') then
                next_state <= decode_instruction;
            end if;
    end case;
end process;

end behavioral;