----------------------------------------------------------------------------------
-- Implementation by Pedro Maat C. Massolino,
-- hereby denoted as "the implementer".
--
-- To the extent possible under law, the implementer has waived all copyright
-- and related or neighboring rights to the source code in this file.
-- http://creativecommons.org/publicdomain/zero/1.0/
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

architecture compact_memory_based_v2 of carmela_state_machine_v128 is

type romtype is array(integer range <>) of std_logic_vector(53 downto 0);

constant rom_state_machine_program : romtype(0 to 2261) := (
--  (0) multiplication_direct_0
-- -- In case of size 1
-- reg_a = a0_X; reg_b = b0_X; reg_acc = 0; o0_X = reg_o; o1_X = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001000001110000100000010001100100000000000011",
--  (1) multiplication_direct_1
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (2) multiplication_direct_2
-- -- Other cases
-- reg_a = a0_X; reg_b = b0_X; reg_acc = 0; o0_X = reg_o; operation : a*b + acc; o0_X = reg_o;
"000010100001001000010000100000010000000100000000000011",
--  (3) multiplication_direct_3
-- -- In case of size 2
-- reg_a = a1_X; reg_b = b0_X; reg_acc = reg_o >> 256; Enable sign a; operation : a*b + acc;
"000000100001001000000000100000100000101000100000100011",
--  (4) multiplication_direct_4
-- reg_a = a0_X; reg_b = b1_X; reg_acc = reg_o; o1_X = reg_o; Enable sign b; operation : a*b + acc;
"000000100001001000010000100000000001001000100100000011",
--  (5) multiplication_direct_5
-- reg_a = a1_X; reg_b = b1_X; reg_acc = reg_o >> 256; o2_X = reg_o; o3_X = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001001001110000100000100000001101000100100011",
--  (6) multiplication_direct_6
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (7) multiplication_direct_7
-- -- Other cases
-- reg_a = a1_X; reg_b = b0_X; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001010000000000100000100000001000100000100011",
--  (8) multiplication_direct_8
-- reg_a = a0_X; reg_b = b1_X; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
"000000100001010000010000100000000000001000100100000011",
--  (9) multiplication_direct_9
-- reg_a = a1_X; reg_b = b1_X; reg_acc = reg_o >> 256; operation : a*b + acc;
"000011100001010000000000100000100000001101000100100011",
--  (10) multiplication_direct_10
-- -- In case of size 3
-- reg_a = a0_X; reg_b = b2_X; reg_acc = reg_o; Enable sign b; operation : a*b + acc;
"000000100001010000000000100000000001001101001000000011",
--  (11) multiplication_direct_11
-- reg_a = a2_X; reg_b = b0_X; reg_acc = reg_o; Enable sign a; o2_X = reg_o; operation : a*b + acc;
"000000100001010000010000100000000000101101000001000011",
--  (12) multiplication_direct_12
-- reg_a = a2_X; reg_b = b1_X; reg_acc = reg_o >> 256; Enable sign a; operation : a*b + acc;
"000000100001010000000000100000100000110001100101000011",
--  (13) multiplication_direct_13
-- reg_a = a1_X; reg_b = b2_X; reg_acc = reg_o; o3_X = reg_o; Enable sign b; operation : a*b + acc;
"000000100001010000010000100000000001010001101000100011",
--  (14) multiplication_direct_14
-- reg_a = a2_X; reg_b = b2_X; reg_acc = reg_o >> 256; o4_X = reg_o; o5_X = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001010001110000100000100001110110001001000011",
--  (15) multiplication_direct_15
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (16) multiplication_direct_16
-- -- Other cases
-- reg_a = a0_0; reg_b = b2_0; reg_acc = reg_o; operation : a*b + acc;
"000000100001011000000000100000000000001101001000000011",
--  (17) multiplication_direct_17
-- reg_a = a2_X; reg_b = b0_X; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
"000000100001011000010000100000000000001101000001000011",
--  (18) multiplication_direct_18
-- reg_a = a2_X; reg_b = b1_X; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001011000000000100000100000010001100101000011",
--  (19) multiplication_direct_19
-- reg_a = a1_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000101000001011000000000100000000000010001101000100011",
--  (20) multiplication_direct_20
-- -- In case of size 4
-- reg_a = a3_X; reg_b = b0_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001011000000000100000000000110001100001100011",
--  (21) multiplication_direct_21
-- reg_a = a0_X; reg_b = b3_X; reg_acc = reg_o; o3_X = reg_o; Enable sign b; operation : a*b + acc;
"000000100001011000010000100000000001010001101100000011",
--  (22) multiplication_direct_22
-- reg_a = a2_X; reg_b = b2_X; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001011000000000100000100000010110001001000011",
--  (23) multiplication_direct_23
-- reg_a = a3_X; reg_b = b1_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001011000000000100000000000110110000101100011",
--  (24) multiplication_direct_24
-- reg_a = a1_X; reg_b = b3_X; reg_acc = reg_o; o4_X = reg_o; Enable sign b; operation : a*b + acc;
"000000100001011000010000100000000001010110001100100011",
--  (25) multiplication_direct_25
-- reg_a = a3_X; reg_b = b2_X; reg_acc = reg_o >> 256; Enable sign a; operation : a*b + acc;
"000000100001011000000000100000100000111010101001100011",
--  (26) multiplication_direct_26
-- reg_a = a2_X; reg_b = b3_X; reg_acc = reg_o; o5_X = reg_o; Enable sign b; operation : a*b + acc;
"000000100001011000010000100000000001011010101101000011",
--  (27) multiplication_direct_27
-- reg_a = a3_X; reg_b = b3_X; reg_acc = reg_o >> 256; o6_X = reg_o; o7_X = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001011001110000100000100001111111001101100011",
--  (28) multiplication_direct_28
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (29) multiplication_direct_29
-- -- Other cases
-- reg_a = a3_X; reg_b = b0_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000010001100001100011",
--  (30) multiplication_direct_30
-- reg_a = a0_X; reg_b = b3_X; reg_acc = reg_o; o3_0 = reg_o; operation : a*b + acc;
"000000100001100000010000100000000000010001101100000011",
--  (31) multiplication_direct_31
-- reg_a = a2_X; reg_b = b2_X; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001100000000000100000100000010110001001000011",
--  (32) multiplication_direct_32
-- reg_a = a3_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000010110000101100011",
--  (33) multiplication_direct_33
-- reg_a = a1_X; reg_b = b3_X; reg_acc = reg_o; o4_0 = reg_o; operation : a*b + acc;
"000111000001100000010000100000000000010110001100100011",
--  (34) multiplication_direct_34
-- -- In case of size 5
-- reg_a = a4_X; reg_b = b0_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001100000000000100000000000110110000010000011",
--  (35) multiplication_direct_35
-- reg_a = a0_X; reg_b = b4_X; reg_acc = reg_o; o4_0 = reg_o; Enable sign b; operation : a*b + acc;
"000000100001100000010000100000000001010110010000000011",
--  (36) multiplication_direct_36
-- reg_a = a3_X; reg_b = b2_X; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001100000000000100000100000011010101001100011",
--  (37) multiplication_direct_37
-- reg_a = a2_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000011010101101000011",
--  (38) multiplication_direct_38
-- reg_a = a4_X; reg_b = b1_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001100000000000100000000000111010100110000011",
--  (39) multiplication_direct_39
-- reg_a = a1_X; reg_b = b4_X; reg_acc = reg_o; o5_X = reg_o; Enable sign b; operation : a*b + acc;
"000000100001100000010000100000000001011010110000100011",
--  (40) multiplication_direct_40
-- reg_a = a3_X; reg_b = b3_X; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001100000000000100000100000011111001101100011",
--  (41) multiplication_direct_41
-- reg_a = a4_X; reg_b = b2_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001100000000000100000000000111111001010000011",
--  (42) multiplication_direct_42
-- reg_a = a2_X; reg_b = b4_X; reg_acc = reg_o; o6_X = reg_o; Enable sign b; operation : a*b + acc;
"000000100001100000010000100000000001011111010001000011",
--  (43) multiplication_direct_43
-- reg_a = a4_X; reg_b = b3_X; reg_acc = reg_o >> 256; Enable sign a; operation : a*b + acc;
"000000100001100000000000100000100000100011101110000011",
--  (44) multiplication_direct_44
-- reg_a = a3_X; reg_b = b4_X; reg_acc = reg_o; o7_X = reg_o; Enable sign b; operation : a*b + acc; Increment base address o;
"000000100001100010010000100000000001000011110001100011",
--  (45) multiplication_direct_45
-- reg_a = a4_X; reg_b = b4_X; reg_acc = reg_o >> 256; o8_X = reg_o; o9_X = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001100001110000100000100001100100010010000011",
--  (46) multiplication_direct_46
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (47) multiplication_direct_47
-- -- Other cases
-- reg_a = a4_X; reg_b = b0_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000010110000010000011",
--  (48) multiplication_direct_48
-- reg_a = a0_X; reg_b = b4_X; reg_acc = reg_o; o4_X = reg_o; operation : a*b + acc;
"000000100001101000010000100000000000010110010000000011",
--  (49) multiplication_direct_49
-- reg_a = a3_X; reg_b = b2_X; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001101000000000100000100000011010101001100011",
--  (50) multiplication_direct_50
-- reg_a = a2_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000011010101101000011",
--  (51) multiplication_direct_51
-- reg_a = a4_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000011010100110000011",
--  (52) multiplication_direct_52
-- reg_a = a1_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"001001100001101000000000100000000000011010110000100011",
--  (53) multiplication_direct_53
-- -- In case of size 6
-- reg_a = a5_X; reg_b = b0_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001101000000000100000000000111010100010100011",
--  (54) multiplication_direct_54
-- reg_a = a0_X; reg_b = b5_X; reg_acc = reg_o; o5_0 = reg_o; Enable sign b; operation : a*b + acc;
"000000100001101000010000100000000001011010110100000011",
--  (55) multiplication_direct_55
-- reg_a = a3_X; reg_b = b3_X; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001101000000000100000100000011111001101100011",
--  (56) multiplication_direct_56
-- reg_a = a2_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000011111010001000011",
--  (57) multiplication_direct_57
-- reg_a = a4_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000011111001010000011",
--  (58) multiplication_direct_58
-- reg_a = a5_X; reg_b = b1_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001101000000000100000000000111111000110100011",
--  (59) multiplication_direct_59
-- reg_a = a1_X; reg_b = b5_X; reg_acc = reg_o; o6_0 = reg_o; Enable sign b; operation : a*b + acc;
"000000100001101000010000100000000001011111010100100011",
--  (60) multiplication_direct_60
-- reg_a = a4_X; reg_b = b3_X; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001101000000000100000100000000011101110000011",
--  (61) multiplication_direct_61
-- reg_a = a3_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000011110001100011",
--  (62) multiplication_direct_62
-- reg_a = a5_X; reg_b = b2_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001101000000000100000000000100011101010100011",
--  (63) multiplication_direct_63
-- reg_a = a2_X; reg_b = b5_X; reg_acc = reg_o; o7_0 = reg_o; Enable sign b; operation : a*b + acc; Increment base address o;
"000000100001101010010000100000000001000011110101000011",
--  (64) multiplication_direct_64
-- reg_a = a4_X; reg_b = b4_X; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001101000000000100000100000000100010010000011",
--  (65) multiplication_direct_65
-- reg_a = a5_X; reg_b = b3_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001101000000000100000000000100100001110100011",
--  (66) multiplication_direct_66
-- reg_a = a3_X; reg_b = b5_X; reg_acc = reg_o; o8_0 = reg_o; Enable sign b; operation : a*b + acc;
"000000100001101000010000100000000001000100010101100011",
--  (67) multiplication_direct_67
-- reg_a = a5_X; reg_b = b4_X; reg_acc = reg_o >> 256; Enable sign a; operation : a*b + acc;
"000000100001101000000000100000100000101000110010100011",
--  (68) multiplication_direct_68
-- reg_a = a4_X; reg_b = b5_X; reg_acc = reg_o; o9_0 = reg_o; Enable sign b; operation : a*b + acc;
"000000100001101000010000100000000001001000110110000011",
--  (69) multiplication_direct_69
-- reg_a = a5_X; reg_b = b5_X; reg_acc = reg_o >> 256; o10_X = reg_o; o11_X = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001101001110000100000100001101101010110100011",
--  (70) multiplication_direct_70
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (71) multiplication_direct_71
-- -- Other cases
-- reg_a = a5_X; reg_b = b0_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000011010100010100011",
--  (72) multiplication_direct_72
-- reg_a = a0_X; reg_b = b5_X; reg_acc = reg_o; o5_0 = reg_o; operation : a*b + acc;
"000000100001110000010000100000000000011010110100000011",
--  (73) multiplication_direct_73
-- reg_a = a3_X; reg_b = b3_X; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001110000000000100000100000011111001101100011",
--  (74) multiplication_direct_74
-- reg_a = a4_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000011111001010000011",
--  (75) multiplication_direct_75
-- reg_a = a2_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000011111010001000011",
--  (76) multiplication_direct_76
-- reg_a = a5_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000011111000110100011",
--  (77) multiplication_direct_77
-- reg_a = a1_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"001100100001110000000000100000000000011111010100100011",
--  (78) multiplication_direct_78
-- -- In case of size 7
-- reg_a = a6_X; reg_b = b0_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001110000000000100000000000111111000011000011",
--  (79) multiplication_direct_79
-- reg_a = a0_X; reg_b = b6_X; reg_acc = reg_o; o6_0 = reg_o; Enable sign b; operation : a*b + acc;
"000000100001110000010000100000000001011111011000000011",
--  (80) multiplication_direct_80
-- reg_a = a4_X; reg_b = b3_X; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001110000000000100000100000000011101110000011",
--  (81) multiplication_direct_81
-- reg_a = a3_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000011110001100011",
--  (82) multiplication_direct_82
-- reg_a = a5_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000011101010100011",
--  (83) multiplication_direct_83
-- reg_a = a2_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000011110101000011",
--  (84) multiplication_direct_84
-- reg_a = a6_X; reg_b = b1_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001110000000000100000000000100011100111000011",
--  (85) multiplication_direct_85
-- reg_a = a1_X; reg_b = b6_X; reg_acc = reg_o; o7_0 = reg_o; Enable sign b; operation : a*b + acc; Increment base address o;
"000000100001110010010000100000000001000011111000100011",
--  (86) multiplication_direct_86
-- reg_a = a4_X; reg_b = b4_X; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001110000000000100000100000000100010010000011",
--  (87) multiplication_direct_87
-- reg_a = a5_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001110100011",
--  (88) multiplication_direct_88
-- reg_a = a3_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010101100011",
--  (89) multiplication_direct_89
-- reg_a = a6_X; reg_b = b2_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001110000000000100000000000100100001011000011",
--  (90) multiplication_direct_90
-- reg_a = a2_X; reg_b = b6_X; reg_acc = reg_o; o8_0 = reg_o; Enable sign b; operation : a*b + acc;
"000000100001110000010000100000000001000100011001000011",
--  (91) multiplication_direct_91
-- reg_a = a5_X; reg_b = b4_X; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001110000000000100000100000001000110010100011",
--  (92) multiplication_direct_92
-- reg_a = a4_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000001000110110000011",
--  (93) multiplication_direct_93
-- reg_a = a6_X; reg_b = b3_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001110000000000100000000000101000101111000011",
--  (94) multiplication_direct_94
-- reg_a = a3_X; reg_b = b6_X; reg_acc = reg_o; o9_0 = reg_o; Enable sign b; operation : a*b + acc;
"000000100001110000010000100000000001001000111001100011",
--  (95) multiplication_direct_95
-- reg_a = a5_X; reg_b = b5_X; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001110000000000100000100000001101010110100011",
--  (96) multiplication_direct_96
-- reg_a = a6_X; reg_b = b4_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001110000000000100000000000101101010011000011",
--  (97) multiplication_direct_97
-- reg_a = a4_X; reg_b = b6_X; reg_acc = reg_o; o10_0 = reg_o; Enable sign b; operation : a*b + acc;
"000000100001110000010000100000000001001101011010000011",
--  (98) multiplication_direct_98
-- reg_a = a6_X; reg_b = b5_X; reg_acc = reg_o >> 256; Enable sign a; operation : a*b + acc;
"000000100001110000000000100000100000110001110111000011",
--  (99) multiplication_direct_99
-- reg_a = a5_X; reg_b = b6_X; reg_acc = reg_o; o11_0 = reg_o; Enable sign b; operation : a*b + acc;
"000000100001110000010000100000000001010001111010100011",
--  (100) multiplication_direct_100
-- reg_a = a6_X; reg_b = b6_X; reg_acc = reg_o >> 256; o12_X = reg_o; o13_X = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001110001110000100000100001110110011011000011",
--  (101) multiplication_direct_101
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (102) multiplication_direct_102
-- -- In case of size 8
-- reg_a = a6_X; reg_b = b0_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000011111000011000011",
--  (103) multiplication_direct_103
-- reg_a = a0_X; reg_b = b6_X; reg_acc = reg_o; o6_0 = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000011111011000000011",
--  (104) multiplication_direct_104
-- reg_a = a4_X; reg_b = b3_X; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001111000000000100000100000000011101110000011",
--  (105) multiplication_direct_105
-- reg_a = a3_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000011110001100011",
--  (106) multiplication_direct_106
-- reg_a = a5_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000011101010100011",
--  (107) multiplication_direct_107
-- reg_a = a2_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000011110101000011",
--  (108) multiplication_direct_108
-- reg_a = a6_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000011100111000011",
--  (109) multiplication_direct_109
-- reg_a = a1_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000011111000100011",
--  (110) multiplication_direct_110
-- reg_a = a7_X; reg_b = b0_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001111000000000100000000000100011100011100011",
--  (111) multiplication_direct_111
-- reg_a = a0_X; reg_b = b7_X; reg_acc = reg_o; o7_0 = reg_o; Enable sign b; operation : a*b + acc; Increment base address o;
"000000100001111010010000100000000001000011111100000011",
--  (112) multiplication_direct_112
-- reg_a = a4_X; reg_b = b4_X; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001111000000000100000100000000100010010000011",
--  (113) multiplication_direct_113
-- reg_a = a5_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001110100011",
--  (114) multiplication_direct_114
-- reg_a = a3_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010101100011",
--  (115) multiplication_direct_115
-- reg_a = a6_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001011000011",
--  (116) multiplication_direct_116
-- reg_a = a2_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011001000011",
--  (117) multiplication_direct_117
-- reg_a = a7_X; reg_b = b1_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001111000000000100000000000100100000111100011",
--  (118) multiplication_direct_118
-- reg_a = a1_X; reg_b = b7_X; reg_acc = reg_o; o8_0 = reg_o; Enable sign b; operation : a*b + acc;
"000000100001111000010000100000000001000100011100100011",
--  (119) multiplication_direct_119
-- reg_a = a5_X; reg_b = b4_X; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001111000000000100000100000001000110010100011",
--  (120) multiplication_direct_120
-- reg_a = a4_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000001000110110000011",
--  (121) multiplication_direct_121
-- reg_a = a6_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000001000101111000011",
--  (122) multiplication_direct_122
-- reg_a = a3_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000001000111001100011",
--  (123) multiplication_direct_123
-- reg_a = a7_X; reg_b = b2_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001111000000000100000000000101000101011100011",
--  (124) multiplication_direct_124
-- reg_a = a2_X; reg_b = b7_X; reg_acc = reg_o; o9_0 = reg_o; Enable sign b; operation : a*b + acc;
"000000100001111000010000100000000001001000111101000011",
--  (125) multiplication_direct_125
-- reg_a = a5_X; reg_b = b5_X; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001111000000000100000100000001101010110100011",
--  (126) multiplication_direct_126
-- reg_a = a6_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000001101010011000011",
--  (127) multiplication_direct_127
-- reg_a = a4_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000001101011010000011",
--  (128) multiplication_direct_128
-- reg_a = a7_X; reg_b = b3_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001111000000000100000000000101101001111100011",
--  (129) multiplication_direct_129
-- reg_a = a3_X; reg_b = b7_X; reg_acc = reg_o; o10_0 = reg_o; Enable sign b; operation : a*b + acc;
"000000100001111000010000100000000001001101011101100011",
--  (130) multiplication_direct_130
-- reg_a = a6_X; reg_b = b5_X; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001111000000000100000100000010001110111000011",
--  (131) multiplication_direct_131
-- reg_a = a5_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000010001111010100011",
--  (132) multiplication_direct_132
-- reg_a = a7_X; reg_b = b4_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001111000000000100000000000110001110011100011",
--  (133) multiplication_direct_133
-- reg_a = a4_X; reg_b = b7_X; reg_acc = reg_o; o11_0 = reg_o; Enable sign b; operation : a*b + acc;
"000000100001111000010000100000000001010001111110000011",
--  (134) multiplication_direct_134
-- reg_a = a6_X; reg_b = b6_X; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001111000000000100000100000010110011011000011",
--  (135) multiplication_direct_135
-- reg_a = a7_X; reg_b = b5_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001111000000000100000000000110110010111100011",
--  (136) multiplication_direct_136
-- reg_a = a5_X; reg_b = b7_X; reg_acc = reg_o; o12_0 = reg_o; Enable sign b; operation : a*b + acc;
"000000100001111000010000100000000001010110011110100011",
--  (137) multiplication_direct_137
-- reg_a = a7_X; reg_b = b6_X; reg_acc = reg_o >> 256; Enable sign a; operation : a*b + acc;
"000000100001111000000000100000100000111010111011100011",
--  (138) multiplication_direct_138
-- reg_a = a6_X; reg_b = b7_X; reg_acc = reg_o; o13_0 = reg_o; Enable sign b; operation : a*b + acc;
"000000100001111000010000100000000001011010111111000011",
--  (139) multiplication_direct_139
-- reg_a = a7_X; reg_b = b7_X; reg_acc = reg_o >> 256; o14_X = reg_o; o15_X = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001111001110000100000100001111111011111100011",
--  (140) multiplication_direct_140
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (141) square_direct_0
-- -- In case of size 1
-- reg_a = a0_X; reg_b = a0_X; reg_acc = 0; o0_X = reg_o; o1_X = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001000001110000100000010001100100000000000011",
--  (142) square_direct_1
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (143) square_direct_2
-- -- In case of sizes 2, 3, 4, 5, 6, 7, 8
-- reg_a = a0_X; reg_b = a0_X; reg_acc = 0; o0_X = reg_o; operation : a*b + acc;
"000010000001001000010000100000010000000100000000000011",
--  (144) square_direct_3
-- -- In case of size 2
-- reg_a = a1_X; reg_b = a0_X; reg_acc = reg_o >> 256; o1_X = reg_o; Enable sign a; operation : 2*a*b + acc;
"000000100001001000010100100000100000101000100000100011",
--  (145) square_direct_4
-- reg_a = a1_X; reg_b = a1_X; reg_acc = reg_o >> 256; o2_X = reg_o; o3_X = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001001001110000100000100001101101000100100011",
--  (146) square_direct_5
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (147) square_direct_6
-- -- Other cases
-- reg_a = a1_X; reg_b = a0_X; reg_acc = reg_o >> 256; o1_X = reg_o; operation : 2*a*b + acc;
"000000100001010000010100100000100000001000100000100011",
--  (148) square_direct_7
-- reg_a = a1_X; reg_b = a1_X; reg_acc = reg_o >> 256; operation : a*b + acc;
"000010100001010000000000100000100000001101000100100011",
--  (149) square_direct_8
-- -- In case of size 3
-- reg_a = a0_X; reg_b = a2_X; reg_acc = reg_o; o2_X = reg_o; Enable sign b; operation : 2*a*b + acc;
"000000100001010000010100100000000001001101001000000011",
--  (150) square_direct_9
-- reg_a = a2_X; reg_b = a1_X; reg_acc = reg_o >> 256; o3_X = reg_o; Enable sign a; operation : 2*a*b + acc;
"000000100001010000010100100000100000110001100101000011",
--  (151) square_direct_10
-- reg_a = a2_X; reg_b = a2_X; reg_acc = reg_o >> 256; o4_X = reg_o; o5_X = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001010001110000100000100001110110001001000011",
--  (152) square_direct_11
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (153) square_direct_12
-- -- Other cases
-- reg_a = a0_X; reg_b = a2_X; reg_acc = reg_o; o2_X = reg_o; operation : 2*a*b + acc;
"000000100001011000010100100000000000001101001000000011",
--  (154) square_direct_13
-- reg_a = a2_X; reg_b = a1_X; reg_acc = reg_o >> 256; operation : 2*a*b + acc;
"000011100001011000000100100000100000010001100101000011",
--  (155) square_direct_14
-- -- In case of size 4
-- reg_a = a3_X; reg_b = a0_X; reg_acc = reg_o; o3_X = reg_o; Enable sign a; operation : 2*a*b + acc;
"000000100001011000010100100000000000110001100001100011",
--  (156) square_direct_15
-- reg_a = a2_X; reg_b = a2_X; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001011000000000100000100000010110001001000011",
--  (157) square_direct_16
-- reg_a = a3_X; reg_b = a1_X; reg_acc = reg_o; o4_X = reg_o; Enable sign a; operation : 2*a*b + acc;
"000000100001011000010100100000000000110110000101100011",
--  (158) square_direct_17
-- reg_a = a3_X; reg_b = a2_X; reg_acc = reg_o >> 256; o5_X = reg_o; Enable sign a; operation : 2*a*b + acc;
"000000100001011000010100100000100000111010101001100011",
--  (159) square_direct_18
-- reg_a = a3_X; reg_b = a3_X; reg_acc = reg_o >> 256; o6_X = reg_o; o7_X = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001011001110000100000100001111111001101100011",
--  (160) square_direct_19
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (161) square_direct_20
-- -- Other cases
-- reg_a = a3_X; reg_b = a0_X; reg_acc = reg_o; o3_X = reg_o; operation : 2*a*b + acc;
"000000100001100000010100100000000000010001100001100011",
--  (162) square_direct_21
-- reg_a = a2_X; reg_b = a2_X; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001100000000000100000100000010110001001000011",
--  (163) square_direct_22
-- reg_a = a3_X; reg_b = a1_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000100100001100000000100100000000000010110000101100011",
--  (164) square_direct_23
-- -- In case of size 5
-- reg_a = a4_X; reg_b = a0_X; reg_acc = reg_o; o4_X = reg_o; Enable sign a; operation : 2*a*b + acc;
"000000100001100000010100100000000000110110000010000011",
--  (165) square_direct_24
-- reg_a = a3_X; reg_b = a2_X; reg_acc = reg_o >> 256; operation : 2*a*b + acc;
"000000100001100000000100100000100000011010101001100011",
--  (166) square_direct_25
-- reg_a = a4_X; reg_b = a1_X; reg_acc = reg_o; o5_X = reg_o; Enable sign a; operation : 2*a*b + acc;
"000000100001100000010100100000000000111010100110000011",
--  (167) square_direct_26
-- reg_a = a3_X; reg_b = a3_X; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001100000000000100000100000011111011011000011",
--  (168) square_direct_27
-- reg_a = a4_X; reg_b = a2_X; reg_acc = reg_o; o6_X = reg_o; Enable sign a; operation : 2*a*b + acc;
"000000100001100000010100100000000000111111001010000011",
--  (169) square_direct_28
-- reg_a = a4_X; reg_b = a3_X; reg_acc = reg_o >> 256; o7_X = reg_o; Enable sign a; operation : 2*a*b + acc; Increase base address o;
"000000100001100010010100100000100000100011101110000011",
--  (170) square_direct_29
-- reg_a = a4_X; reg_b = a4_X; reg_acc = reg_o >> 256; o8_X = reg_o; o9_X = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001100001110000100000100001100100010010000011",
--  (171) square_direct_30
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (172) square_direct_31
-- -- Other cases
-- reg_a = a4_X; reg_b = a0_X; reg_acc = reg_o; o4_X = reg_o; operation : 2*a*b + acc;
"000000100001101000010100100000000000010110000010000011",
--  (173) square_direct_32
-- reg_a = a3_X; reg_b = a2_X; reg_acc = reg_o >> 256; operation : 2*a*b + acc;
"000000100001101000000100100000100000010110001001100011",
--  (174) square_direct_33
-- reg_a = a4_X; reg_b = a1_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000110000001101000000100100000000000011010100110000011",
--  (175) square_direct_34
-- -- In case of size 6
-- reg_a = a5_X; reg_b = a0_X; reg_acc = reg_o; o5_X = reg_o; Enable sign a; operation : 2*a*b + acc;
"000000100001101000010100100000000000111010100010100011",
--  (176) square_direct_35
-- reg_a = a3_X; reg_b = a3_X; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001101000000000100000100000011111001101100011",
--  (177) square_direct_36
-- reg_a = a4_X; reg_b = a2_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001101000000100100000000000011111001010000011",
--  (178) square_direct_37
-- reg_a = a5_X; reg_b = a1_X; reg_acc = reg_o; o6_X = reg_o; Enable sign a; operation : 2*a*b + acc;
"000000100001101000010100100000000000111011000110100011",
--  (179) square_direct_38
-- reg_a = a4_X; reg_b = a3_X; reg_acc = reg_o >> 256; operation : 2*a*b + acc;
"000000100001101000000100100000100000000011101110000011",
--  (180) square_direct_39
-- reg_a = a5_X; reg_b = a2_X; reg_acc = reg_o; o7_X = reg_o; Enable sign a; operation : 2*a*b + acc; Increase base address o;
"000000100001101010010100100000000000100011101010100011",
--  (181) square_direct_40
-- reg_a = a4_X; reg_b = a4_X; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001101000000000100000100000000100010010000011",
--  (182) square_direct_41
-- reg_a = a5_X; reg_b = a3_X; reg_acc = reg_o; o8_X = reg_o; Enable sign a; operation : 2*a*b + acc;
"000000100001101000010100100000000000100100001110100011",
--  (183) square_direct_42
-- reg_a = a5_X; reg_b = a4_X; reg_acc = reg_o >> 256; o9_X = reg_o; Enable sign a; operation : 2*a*b + acc;
"000000100001101000010100100000100000101000110010100011",
--  (184) square_direct_43
-- reg_a = a5_X; reg_b = a5_X; reg_acc = reg_o >> 256; o10_X = reg_o; o11_X = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001101001110000100000100001101101010110100011",
--  (185) square_direct_44
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (186) square_direct_45
-- -- Other cases
-- reg_a = a5_X; reg_b = a0_X; reg_acc = reg_o; o5_X = reg_o; operation : 2*a*b + acc;
"000000100001110000010100100000000000011010100010100011",
--  (187) square_direct_46
-- reg_a = a3_X; reg_b = a3_X; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001110000000000100000100000011111001101100011",
--  (188) square_direct_47
-- reg_a = a4_X; reg_b = a2_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001110000000100100000000000011111001010000011",
--  (189) square_direct_48
-- reg_a = a5_X; reg_b = a1_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000111100001110000000100100000000000011111000110100011",
--  (190) square_direct_49
-- -- In case of size 7
-- reg_a = a6_X; reg_b = a0_X; reg_acc = reg_o; o6_X = reg_o; Enable sign a; operation : 2*a*b + acc;
"000000100001110000010100100000000000111111000011000011",
--  (191) square_direct_50
-- reg_a = a4_X; reg_b = a3_X; reg_acc = reg_o >> 256; operation : 2*a*b + acc;
"000000100001110000000100100000100000000011101110000011",
--  (192) square_direct_51
-- reg_a = a5_X; reg_b = a2_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001110000000100100000000000000011101010100011",
--  (193) square_direct_52
-- reg_a = a6_X; reg_b = a1_X; reg_acc = reg_o; o7_X = reg_o; Enable sign a; operation : 2*a*b + acc; Increase base address o;
"000000100001110010010100100000000000100011100111000011",
--  (194) square_direct_53
-- reg_a = a4_X; reg_b = a4_X; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001110000000000100000100000000100010010000011",
--  (195) square_direct_54
-- reg_a = a5_X; reg_b = a3_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001110000000100100000000000000100001110100011",
--  (196) square_direct_55
-- reg_a = a6_X; reg_b = a2_X; reg_acc = reg_o; o8_X = reg_o; Enable sign a; operation : 2*a*b + acc;
"000000100001110000010100100000000000100100001011000011",
--  (197) square_direct_56
-- reg_a = a5_X; reg_b = a4_X; reg_acc = reg_o >> 256; operation : 2*a*b + acc;
"000000100001110000000100100000100000001000110010100011",
--  (198) square_direct_57
-- reg_a = a6_X; reg_b = a3_X; reg_acc = reg_o; o9_X = reg_o; Enable sign a; operation : 2*a*b + acc;
"000000100001110000010100100000000000101000101111000011",
--  (199) square_direct_58
-- reg_a = a5_X; reg_b = a5_X; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001110000000000100000100000001101010110100011",
--  (200) square_direct_59
-- reg_a = a6_X; reg_b = a4_X; reg_acc = reg_o; o10_X = reg_o; Enable sign a; operation : 2*a*b + acc;
"000000100001110000010100100000000000101101010011000011",
--  (201) square_direct_60
-- reg_a = a6_X; reg_b = a5_X; reg_acc = reg_o >> 256; o11_X = reg_o; Enable sign a; operation : 2*a*b + acc;
"000000100001110000010100100000100000110001110111000011",
--  (202) square_direct_61
-- reg_a = a6_X; reg_b = a6_X; reg_acc = reg_o >> 256; o12_X = reg_o; o13_X = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001110001110000100000100001110110011011000011",
--  (203) square_direct_62
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (204) square_direct_63
-- -- In case of size 8
-- reg_a = a6_X; reg_b = a0_X; reg_acc = reg_o; o6_X = reg_o; operation : 2*a*b + acc;
"000000100001111000010100100000000000011111000011000011",
--  (205) square_direct_64
-- reg_a = a4_X; reg_b = a3_X; reg_acc = reg_o >> 256; operation : 2*a*b + acc;
"000000100001111000000100100000100000000011101110000011",
--  (206) square_direct_65
-- reg_a = a5_X; reg_b = a2_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001111000000100100000000000000011101010100011",
--  (207) square_direct_66
-- reg_a = a6_X; reg_b = a1_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001111000000100100000000000000011100111000011",
--  (208) square_direct_67
-- reg_a = a7_X; reg_b = a0_X; reg_acc = reg_o; o7_X = reg_o; Enable sign a; operation : 2*a*b + acc; Increase base address o;
"000000100001111010010100100000000000100011100011100011",
--  (209) square_direct_68
-- reg_a = a4_X; reg_b = a4_X; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001111000000000100000100000000100010010000011",
--  (210) square_direct_69
-- reg_a = a5_X; reg_b = a3_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001111000000100100000000000000100001110100011",
--  (211) square_direct_70
-- reg_a = a6_X; reg_b = a2_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001111000000100100000000000000100001011000011",
--  (212) square_direct_71
-- reg_a = a7_X; reg_b = a1_X; reg_acc = reg_o; o8_X = reg_o; Enable sign a; operation : 2*a*b + acc;
"000000100001111000010100100000000000100100000111100011",
--  (213) square_direct_72
-- reg_a = a5_X; reg_b = a4_X; reg_acc = reg_o >> 256; operation : 2*a*b + acc;
"000000100001111000000100100000100000001000110010100011",
--  (214) square_direct_73
-- reg_a = a6_X; reg_b = a3_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001111000000100100000000000001000101111000011",
--  (215) square_direct_74
-- reg_a = a7_X; reg_b = a2_X; reg_acc = reg_o; o9_X = reg_o; Enable sign a; operation : 2*a*b + acc;
"000000100001111000010100100000000000101000101011100011",
--  (216) square_direct_75
-- reg_a = a5_X; reg_b = a5_X; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001111000000000100000100000001101010110100011",
--  (217) square_direct_76
-- reg_a = a6_X; reg_b = a4_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001111000000100100000000000001101010011000011",
--  (218) square_direct_77
-- reg_a = a7_X; reg_b = a3_X; reg_acc = reg_o; o10_X = reg_o; Enable sign a; operation : 2*a*b + acc;
"000000100001111000010100100000000000101101001111100011",
--  (219) square_direct_78
-- reg_a = a6_X; reg_b = a5_X; reg_acc = reg_o >> 256; operation : 2*a*b + acc;
"000000100001111000000100100000100000010001110111000011",
--  (220) square_direct_79
-- reg_a = a7_X; reg_b = a4_X; reg_acc = reg_o; o11_X = reg_o; Enable sign a; operation : 2*a*b + acc;
"000000100001111000010100100000000000110001110011100011",
--  (221) square_direct_80
-- reg_a = a6_X; reg_b = a6_X; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001111000000000100000100000010110011011000011",
--  (222) square_direct_81
-- reg_a = a7_X; reg_b = a5_X; reg_acc = reg_o; o12_X = reg_o; Enable sign a; operation : 2*a*b + acc;
"000000100001111000010100100000000000110110010111100011",
--  (223) square_direct_82
-- reg_a = a7_X; reg_b = a6_X; reg_acc = reg_o >> 256; o13_X = reg_o; Enable sign a; operation : 2*a*b + acc;
"000000100001111000010100100000100000111010111011100011",
--  (224) square_direct_83
-- reg_a = a7_X; reg_b = a7_X; reg_acc = reg_o >> 256; o14_X = reg_o; o15_X = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001111001110000100000100001111111011111100011",
--  (225) square_direct_84
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (226) multiplication_with_reduction_0
-- -- In case of size 1
-- reg_a = a0_X; reg_b = b0_X; reg_acc = 0; Enable sign a,b; operation : a*b + acc;
"000000100001000000000000100000010001100100000000000011",
--  (227) multiplication_with_reduction_1
-- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o0_X = reg_y; operation : keep accumulator;
"000000100001000000011000110000000100000100000000011011",
--  (228) multiplication_with_reduction_2
-- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
"000000100001000000000000100000000010000100000000010011",
--  (229) multiplication_with_reduction_3
-- reg_a = 0; reg_b = 0; reg_acc = reg_o >> 256; o0_X = reg_o; operation : a*b + acc;
"000000100001000000010000100000101110000100000000000011",
--  (230) multiplication_with_reduction_4
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (231) multiplication_with_reduction_5
-- -- In case of sizes 2, 3, 4, 5, 6, 7, 8
-- reg_a = a0_X; reg_b = b0_X; reg_acc = 0; operation : a*b + acc;
"000000100001001000000000100000010000000100000000000011",
--  (232) multiplication_with_reduction_6
-- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o0_X = reg_y; operation : keep accumulator;
"000000100001001000011000110000000100000100000000011011",
--  (233) multiplication_with_reduction_7
-- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
"000000100001001000000000100000000010000100000000010011",
--  (234) multiplication_with_reduction_8
--reg_a = o0_X; reg_b = prime1; reg_acc = reg_o >> 256; operation : a*b + acc;
"000100000001001000000000100000100000000100000100010111",
--  (235) multiplication_with_reduction_9
-- -- In case of size 2
-- reg_a = a0_X; reg_b = b1_X; reg_acc = reg_o; Enable sign b; operation : a*b + acc;
"000000100001001000000000100000000001000100000100000011",
--  (236) multiplication_with_reduction_10
-- reg_a = a1_X; reg_b = b0_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001001000000000100000000000100100000000100011",
--  (237) multiplication_with_reduction_11
-- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o1_X = reg_y; operation : keep accumulator;
"000000100001001000011000110000000100001000100000011011",
--  (238) multiplication_with_reduction_12
-- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
"000000100001001000000000100000000010000100000000010011",
--  (239) multiplication_with_reduction_13
-- reg_a = a1_X; reg_b = b1_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001001000000000100000100001100100000100100011",
--  (240) multiplication_with_reduction_14
-- reg_a = o1_X; reg_b = prime1; reg_acc = reg_o; o0_X = reg_o; o1_X = reg_o >> 256; operation : a*b + acc;
"000000100001001001110000100000000000000100000100110111",
--  (241) multiplication_with_reduction_15
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (242) multiplication_with_reduction_16
-- -- Other cases
-- reg_a = a0_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001010000000000100000000000000100000100000011",
--  (243) multiplication_with_reduction_17
-- reg_a = a1_X; reg_b = b0_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001010000000000100000000000000100000000100011",
--  (244) multiplication_with_reduction_18
-- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o1_X = reg_y; operation : keep accumulator;
"000000100001010000011000110000000100001000100000011011",
--  (245) multiplication_with_reduction_19
-- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
"000000100001010000000000100000000010000100000000010011",
--  (246) multiplication_with_reduction_20
-- reg_a = o0_X; reg_b = prime2; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001010000000000100000100000000100001000010111",
--  (247) multiplication_with_reduction_21
-- reg_a = a1_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001010000000000100000000000000100000100100011",
--  (248) multiplication_with_reduction_22
-- reg_a = o1_X; reg_b = prime1; reg_acc = reg_o; operation : a*b + acc;
"000110000001010000000000100000000000000100000100110111",
--  (249) multiplication_with_reduction_23
-- -- In case of size 3
-- reg_a = a0_X; reg_b = b2_X; reg_acc = reg_o; Enable sign b; operation : a*b + acc;
"000000100001010000000000100000000001000100001000000011",
--  (250) multiplication_with_reduction_24
-- reg_a = a2_X; reg_b = b0_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001010000000000100000000000100100000001000011",
--  (251) multiplication_with_reduction_25
-- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o2_X = reg_y; operation : keep accumulator;
"000000100001010000011000110000000100001101000000011011",
--  (252) multiplication_with_reduction_26
-- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
"000000100001010000000000100000000010000100000000010011",
--  (253) multiplication_with_reduction_27
-- reg_a = a1_X; reg_b = b2_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001010000000000100000100001000100001000100011",
--  (254) multiplication_with_reduction_28
-- reg_a = o1_X; reg_b = prime2; reg_acc = reg_o; operation : a*b + acc;
"000000100001010000000000100000000000000100001000110111",
--  (255) multiplication_with_reduction_29
-- reg_a = a2_X; reg_b = b1_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001010000000000100000000000100100000101000011",
--  (256) multiplication_with_reduction_30
-- reg_a = o2_X; reg_b = prime1; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
"000000100001010000010000100000000000000100000101010111",
--  (257) multiplication_with_reduction_31
-- reg_a = a2_X; reg_b = b2_X; reg_acc = reg_o >> 256; Enable sign a, b; operation : a*b + acc;
"000000100001010000000000100000100001100100001001000011",
--  (258) multiplication_with_reduction_32
-- reg_a = o2_X; reg_b = prime2; reg_acc = reg_o; o1_X = reg_o; o2_X = reg_o >> 256; operation : a*b + acc;
"000000100001010001110000100000000000001000101001010111",
--  (259) multiplication_with_reduction_33
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (260) multiplication_with_reduction_34
-- -- Other cases
-- reg_a = a0_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001011000000000100000000000000100001000000011",
--  (261) multiplication_with_reduction_35
-- reg_a = a2_X; reg_b = b0_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001011000000000100000000000000100000001000011",
--  (262) multiplication_with_reduction_36
-- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o2_X = reg_y; operation : keep accumulator;
"000000100001011000011000110000000100001101000000011011",
--  (263) multiplication_with_reduction_37
-- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
"000000100001011000000000100000000010000100000000010011",
--  (264) multiplication_with_reduction_38
-- reg_a = o0_X; reg_b = prime3; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001011000000000100000100000000100001100010111",
--  (265) multiplication_with_reduction_39
-- reg_a = a1_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001011000000000100000000000000100001000100011",
--  (266) multiplication_with_reduction_40
-- reg_a = o1_X; reg_b = prime2; reg_acc = reg_o; operation : a*b + acc;
"000000100001011000000000100000000000000100001000110111",
--  (267) multiplication_with_reduction_41
-- reg_a = a2_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001011000000000100000000000000100000101000011",
--  (268) multiplication_with_reduction_42
-- reg_a = o2_X; reg_b = prime1; reg_acc = reg_o; operation : a*b + acc;
"001001000001011000000000100000000000000100000101010111",
--  (269) multiplication_with_reduction_43
-- -- In case of size 4
-- reg_a = a0_X; reg_b = b3_X; reg_acc = reg_o; Enable sign b; operation : a*b + acc;
"000000100001011000000000100000000001000100001100000011",
--  (270) multiplication_with_reduction_44
-- reg_a = a3_X; reg_b = b0_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001011000000000100000000000100100000001100011",
--  (271) multiplication_with_reduction_45
-- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o3_X = reg_y; operation : keep accumulator;
"000000100001011000011000110000000100000001100000011011",
--  (272) multiplication_with_reduction_46
-- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
"000000100001011000000000100000000010000100000000010011",
--  (273) multiplication_with_reduction_47
-- reg_a = a1_X; reg_b = b3_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001011000000000100000100001000100001100100011",
--  (274) multiplication_with_reduction_48
-- reg_a = o1_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
"000000100001011000000000100000000000000100001100110111",
--  (275) multiplication_with_reduction_49
-- reg_a = a2_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001011000000000100000000000000100001001000011",
--  (276) multiplication_with_reduction_50
-- reg_a = o2_X; reg_b = prime2; reg_acc = reg_o; operation : a*b + acc;
"000000100001011000000000100000000000000100001001010111",
--  (277) multiplication_with_reduction_51
-- reg_a = a3_X; reg_b = b1_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001011000000000100000000000100100000101100011",
--  (278) multiplication_with_reduction_52
-- reg_a = o3_X; reg_b = prime1; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
"000000100001011000010000100000000000000100000101110111",
--  (279) multiplication_with_reduction_53
-- reg_a = a2_X; reg_b = b3_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001011000000000100000100001000100001101000011",
--  (280) multiplication_with_reduction_54
-- reg_a = o2_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
"000000100001011000000000100000000000000100001101010111",
--  (281) multiplication_with_reduction_55
-- reg_a = a3_X; reg_b = b2_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001011000000000100000000000100100001001100011",
--  (282) multiplication_with_reduction_56
-- reg_a = o3_X; reg_b = prime2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
"000000100001011000010000100000000000001000101001110111",
--  (283) multiplication_with_reduction_57
-- reg_a = a3_X; reg_b = b3_X; reg_acc = reg_o >> 256; Enable sign a, b; operation : a*b + acc;
"000000100001011000000000100000100001100100001101100011",
--  (284) multiplication_with_reduction_58
-- reg_a = o3_X; reg_b = prime3; reg_acc = reg_o; o2_X = reg_o; o3_0 = reg_o >> 256; operation : a*b + acc;
"000000100001011001110000100000000000001101001101110111",
--  (285) multiplication_with_reduction_59
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (286) multiplication_with_reduction_60
-- -- Other cases
-- reg_a = a0_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001100000011",
--  (287) multiplication_with_reduction_61
-- reg_a = a3_X; reg_b = b0_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100000001100011",
--  (288) multiplication_with_reduction_62
-- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o3_X = reg_y; operation : keep accumulator;
"000000100001100000011000110000000100010001100000011011",
--  (289) multiplication_with_reduction_63
-- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000010000100000000010011",
--  (290) multiplication_with_reduction_64
-- reg_a = o0_X; reg_b = prime4; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001100000000000100000100000000100010000010111",
--  (291) multiplication_with_reduction_65
-- reg_a = a1_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001100100011",
--  (292) multiplication_with_reduction_66
-- reg_a = o1_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001100110111",
--  (293) multiplication_with_reduction_67
-- reg_a = a2_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001001000011",
--  (294) multiplication_with_reduction_68
-- reg_a = o2_X; reg_b = prime2; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001001010111",
--  (295) multiplication_with_reduction_69
-- reg_a = a3_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100000101100011",
--  (296) multiplication_with_reduction_70
-- reg_a = o3_X; reg_b = prime1; reg_acc = reg_o; operation : a*b + acc;
"001101000001100000000000100000000000000100000101110111",
--  (297) multiplication_with_reduction_71
-- -- In case of size 5
-- reg_a = a0_X; reg_b = b4_X; reg_acc = reg_o; Enable sign b; operation : a*b + acc;
"000000100001100000000000100000000001000100010000000011",
--  (298) multiplication_with_reduction_72
-- reg_a = a4_X; reg_b = b0_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001100000000000100000000000100100000010000011",
--  (299) multiplication_with_reduction_73
-- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o4_X = reg_y; operation : keep accumulator;
"000000100001100000011000110000000100010110000000011011",
--  (300) multiplication_with_reduction_74
-- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000010000100000000010011",
--  (301) multiplication_with_reduction_75
-- reg_a = a1_X; reg_b = b4_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001100000000000100000100001000100010000100011",
--  (302) multiplication_with_reduction_76
-- reg_a = o1_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100010000110111",
--  (303) multiplication_with_reduction_77
-- reg_a = a2_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001101000011",
--  (304) multiplication_with_reduction_78
-- reg_a = o2_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001101010111",
--  (305) multiplication_with_reduction_79
-- reg_a = a3_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001001100011",
--  (306) multiplication_with_reduction_80
-- reg_a = o3_X; reg_b = prime2; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001001110111",
--  (307) multiplication_with_reduction_81
-- reg_a = a4_X; reg_b = b1_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001100000000000100000000000100100000110000011",
--  (308) multiplication_with_reduction_82
-- reg_a = o4_X; reg_b = prime1; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
"000000100001100000010000100000000000000100000110010111",
--  (309) multiplication_with_reduction_83
-- reg_a = a2_X; reg_b = b4_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001100000000000100000100001000100010001000011",
--  (310) multiplication_with_reduction_84
-- reg_a = o2_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100010001010111",
--  (311) multiplication_with_reduction_85
-- reg_a = a3_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001101100011",
--  (312) multiplication_with_reduction_86
-- reg_a = o3_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001101110111",
--  (313) multiplication_with_reduction_87
-- reg_a = a4_X; reg_b = b2_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001100000000000100000000000100100001010000011",
--  (314) multiplication_with_reduction_88
-- reg_a = o4_X; reg_b = prime2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
"000000100001100000010000100000000000001000101010010111",
--  (315) multiplication_with_reduction_89
-- reg_a = a3_X; reg_b = b4_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001100000000000100000100001000100010001100011",
--  (316) multiplication_with_reduction_90
-- reg_a = o3_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100010001110111",
--  (317) multiplication_with_reduction_91
-- reg_a = a4_X; reg_b = b3_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001100000000000100000000000100100001110000011",
--  (318) multiplication_with_reduction_92
-- reg_a = o4_X; reg_b = prime3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
"000000100001100000010000100000000000001101001110010111",
--  (319) multiplication_with_reduction_93
-- reg_a = a4_X; reg_b = b4_X; reg_acc = reg_o >> 256; Enable sign a, b; operation : a*b + acc;
"000000100001100000000000100000100001100100010010000011",
--  (320) multiplication_with_reduction_94
-- reg_a = o4_X; reg_b = prime4; reg_acc = reg_o; o3_X = reg_o; o4_0 = reg_o >> 256; operation : a*b + acc;
"000000100001100001110000100000000000010001110010010111",
--  (321) multiplication_with_reduction_95
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (322) multiplication_with_reduction_96
-- -- Other cases
-- reg_a = a0_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010000000011",
--  (323) multiplication_with_reduction_97
-- reg_a = a4_X; reg_b = b0_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100000010000011",
--  (324) multiplication_with_reduction_98
-- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o4_X = reg_y; operation : keep accumulator;
"000000100001101000011000110000000100010110000000011011",
--  (325) multiplication_with_reduction_99
-- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000010000100000000010011",
--  (326) multiplication_with_reduction_100
-- reg_a = o0_X; reg_b = prime5; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001101000000000100000100000000100010100010111",
--  (327) multiplication_with_reduction_101
-- reg_a = a1_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010000100011",
--  (328) multiplication_with_reduction_102
-- reg_a = o1_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010000110111",
--  (329) multiplication_with_reduction_103
-- reg_a = a2_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001101000011",
--  (330) multiplication_with_reduction_104
-- reg_a = o2_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001101010111",
--  (331) multiplication_with_reduction_105
-- reg_a = a3_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001001100011",
--  (332) multiplication_with_reduction_106
-- reg_a = o3_X; reg_b = prime2; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001001110111",
--  (333) multiplication_with_reduction_107
-- reg_a = a4_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100000110000011",
--  (334) multiplication_with_reduction_108
-- reg_a = o4_X; reg_b = prime1; reg_acc = reg_o; operation : a*b + acc;
"010010000001101000000000100000000000000100000110010111",
--  (335) multiplication_with_reduction_109
-- -- In case of size 6
-- reg_a = a0_X; reg_b = b5_X; reg_acc = reg_o; Enable sign b; operation : a*b + acc;
"000000100001101000000000100000000001000100010100000011",
--  (336) multiplication_with_reduction_110
-- reg_a = a5_X; reg_b = b0_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001101000000000100000000000100100000010100011",
--  (337) multiplication_with_reduction_111
-- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o5_X = reg_y; operation : keep accumulator;
"000000100001101000011000110000000100011010100000011011",
--  (338) multiplication_with_reduction_112
-- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000010000100000000010011",
--  (339) multiplication_with_reduction_113
-- reg_a = a1_X; reg_b = b5_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001101000000000100000100001000100010100100011",
--  (340) multiplication_with_reduction_114
-- reg_a = o1_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010100110111",
--  (341) multiplication_with_reduction_115
-- reg_a = a2_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010001000011",
--  (342) multiplication_with_reduction_116
-- reg_a = o2_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010001010111",
--  (343) multiplication_with_reduction_117
-- reg_a = a3_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001101100011",
--  (344) multiplication_with_reduction_118
-- reg_a = o3_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001101110111",
--  (345) multiplication_with_reduction_119
-- reg_a = a4_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001010000011",
--  (346) multiplication_with_reduction_120
-- reg_a = o4_X; reg_b = prime2; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001010010111",
--  (347) multiplication_with_reduction_121
-- reg_a = a5_X; reg_b = b1_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001101000000000100000000000100100000110100011",
--  (348) multiplication_with_reduction_122
-- reg_a = o5_X; reg_b = prime1; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
"000000100001101000010000100000000000000100000110110111",
--  (349) multiplication_with_reduction_123
-- reg_a = a2_X; reg_b = b5_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001101000000000100000100001000100010101000011",
--  (350) multiplication_with_reduction_124
-- reg_a = o2_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010101010111",
--  (351) multiplication_with_reduction_125
-- reg_a = a3_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010001100011",
--  (352) multiplication_with_reduction_126
-- reg_a = o3_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010001110111",
--  (353) multiplication_with_reduction_127
-- reg_a = a4_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001110000011",
--  (354) multiplication_with_reduction_128
-- reg_a = o4_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001110010111",
--  (355) multiplication_with_reduction_129
-- reg_a = a5_X; reg_b = b2_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001101000000000100000000000100100001010100011",
--  (356) multiplication_with_reduction_130
-- reg_a = o5_X; reg_b = prime2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
"000000100001101000010000100000000000001000101010110111",
--  (357) multiplication_with_reduction_131
-- reg_a = a3_X; reg_b = b5_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001101000000000100000100001000100010101100011",
--  (358) multiplication_with_reduction_132
-- reg_a = o3_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010101110111",
--  (359) multiplication_with_reduction_133
-- reg_a = a4_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010010000011",
--  (360) multiplication_with_reduction_134
-- reg_a = o4_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010010010111",
--  (361) multiplication_with_reduction_135
-- reg_a = a5_X; reg_b = b3_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001101000000000100000000000100100001110100011",
--  (362) multiplication_with_reduction_136
-- reg_a = o5_X; reg_b = prime3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
"000000100001101000010000100000000000001101001110110111",
--  (363) multiplication_with_reduction_137
-- reg_a = a4_X; reg_b = b5_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001101000000000100000100001000100010110000011",
--  (364) multiplication_with_reduction_138
-- reg_a = o4_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010110010111",
--  (365) multiplication_with_reduction_139
-- reg_a = a5_X; reg_b = b4_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001101000000000100000000000100100010010100011",
--  (366) multiplication_with_reduction_140
-- reg_a = o5_X; reg_b = prime4; reg_acc = reg_o; o3_X = reg_o; operation : a*b + acc;
"000000100001101000010000100000000000010001110010110111",
--  (367) multiplication_with_reduction_141
-- reg_a = a5_X; reg_b = b5_X; reg_acc = reg_o >> 256; Enable sign a, b; operation : a*b + acc;
"000000100001101000000000100000100001100100010110100011",
--  (368) multiplication_with_reduction_142
-- reg_a = o5_X; reg_b = prime5; reg_acc = reg_o; o4_X = reg_o; o5_0 = reg_o >> 256; operation : a*b + acc;
"000000100001101001110000100000000000010110010110110111",
--  (369) multiplication_with_reduction_143
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (370) multiplication_with_reduction_144
-- -- Other cases
-- reg_a = a0_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010100000011",
--  (371) multiplication_with_reduction_145
-- reg_a = a5_X; reg_b = b0_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100000010100011",
--  (372) multiplication_with_reduction_146
-- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o5_X = reg_y; operation : keep accumulator;
"000000100001110000011000110000000100011010100000011011",
--  (373) multiplication_with_reduction_147
-- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000010000100000000010011",
--  (374) multiplication_with_reduction_148
-- reg_a = o0_X; reg_b = prime6; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001110000000000100000100000000100011000010111",
--  (375) multiplication_with_reduction_149
-- reg_a = a1_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010100100011",
--  (376) multiplication_with_reduction_150
-- reg_a = o1_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010100110111",
--  (377) multiplication_with_reduction_151
-- reg_a = a2_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010001000011",
--  (378) multiplication_with_reduction_152
-- reg_a = o2_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010001010111",
--  (379) multiplication_with_reduction_153
-- reg_a = a3_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001101100011",
--  (380) multiplication_with_reduction_154
-- reg_a = o3_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001101110111",
--  (381) multiplication_with_reduction_155
-- reg_a = a4_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001010000011",
--  (382) multiplication_with_reduction_156
-- reg_a = o4_X; reg_b = prime2; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001010010111",
--  (383) multiplication_with_reduction_157
-- reg_a = a5_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100000110100011",
--  (384) multiplication_with_reduction_158
-- reg_a = o5_X; reg_b = prime1; reg_acc = reg_o; operation : a*b + acc;
"011000000001110000000000100000000000000100000110110111",
--  (385) multiplication_with_reduction_159
-- -- In case of size 7
-- reg_a = a0_X; reg_b = b6_X; reg_acc = reg_o; Enable sign b; operation : a*b + acc;
"000000100001110000000000100000000001000100011000000011",
--  (386) multiplication_with_reduction_160
-- reg_a = a6_X; reg_b = b0_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001110000000000100000000000100100000011000011",
--  (387) multiplication_with_reduction_161
-- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o6_X = reg_y; operation : keep accumulator;
"000000100001110000011000110000000100011111000000011011",
--  (388) multiplication_with_reduction_162
-- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000010000100000000010011",
--  (389) multiplication_with_reduction_163
-- reg_a = a1_X; reg_b = b6_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001110000000000100000100001000100011000100011",
--  (390) multiplication_with_reduction_164
-- reg_a = o1_X; reg_b = prime6; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100011000110111",
--  (391) multiplication_with_reduction_165
-- reg_a = a2_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010101000011",
--  (392) multiplication_with_reduction_166
-- reg_a = o2_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010101010111",
--  (393) multiplication_with_reduction_167
-- reg_a = a3_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010001100011",
--  (394) multiplication_with_reduction_168
-- reg_a = o3_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010001110111",
--  (395) multiplication_with_reduction_169
-- reg_a = a4_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001110000011",
--  (396) multiplication_with_reduction_170
-- reg_a = o4_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001110010111",
--  (397) multiplication_with_reduction_171
-- reg_a = a5_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001010100011",
--  (398) multiplication_with_reduction_172
-- reg_a = o5_X; reg_b = prime2; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001010110111",
--  (399) multiplication_with_reduction_173
-- reg_a = a6_X; reg_b = b1_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001110000000000100000000000100100000111000011",
--  (400) multiplication_with_reduction_174
-- reg_a = o6_X; reg_b = prime1; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
"000000100001110000010000100000000000000100000111010111",
--  (401) multiplication_with_reduction_175
-- reg_a = a2_X; reg_b = b6_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001110000000000100000100001000100011001000011",
--  (402) multiplication_with_reduction_176
-- reg_a = o2_X; reg_b = prime6; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100011001010111",
--  (403) multiplication_with_reduction_177
-- reg_a = a3_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010101100011",
--  (404) multiplication_with_reduction_178
-- reg_a = o3_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010101110111",
--  (405) multiplication_with_reduction_179
-- reg_a = a4_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010010000011",
--  (406) multiplication_with_reduction_180
-- reg_a = o4_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010010010111",
--  (407) multiplication_with_reduction_181
-- reg_a = a5_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001110100011",
--  (408) multiplication_with_reduction_182
-- reg_a = o5_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001110110111",
--  (409) multiplication_with_reduction_183
-- reg_a = a6_X; reg_b = b2_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001110000000000100000000000100100001011000011",
--  (410) multiplication_with_reduction_184
-- reg_a = o6_X; reg_b = prime2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
"000000100001110000010000100000000000001000101011010111",
--  (411) multiplication_with_reduction_185
-- reg_a = a3_X; reg_b = b6_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001110000000000100000100001000100011001100011",
--  (412) multiplication_with_reduction_186
-- reg_a = o3_X; reg_b = prime6; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100011001110111",
--  (413) multiplication_with_reduction_187
-- reg_a = a4_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010110000011",
--  (414) multiplication_with_reduction_188
-- reg_a = o4_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010110010111",
--  (415) multiplication_with_reduction_189
-- reg_a = a5_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010010100011",
--  (416) multiplication_with_reduction_190
-- reg_a = o5_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010010110111",
--  (417) multiplication_with_reduction_191
-- reg_a = a6_X; reg_b = b3_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001110000000000100000000000100100001111000011",
--  (418) multiplication_with_reduction_192
-- reg_a = o6_X; reg_b = prime3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
"000000100001110000010000100000000000001101001111010111",
--  (419) multiplication_with_reduction_193
-- reg_a = a4_X; reg_b = b6_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001110000000000100000100001000100011010000011",
--  (420) multiplication_with_reduction_194
-- reg_a = o4_X; reg_b = prime6; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100011010010111",
--  (421) multiplication_with_reduction_195
-- reg_a = a5_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010110100011",
--  (422) multiplication_with_reduction_196
-- reg_a = o5_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010110110111",
--  (423) multiplication_with_reduction_197
-- reg_a = a6_X; reg_b = b4_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001110000000000100000000000100100010011000011",
--  (424) multiplication_with_reduction_198
-- reg_a = o6_X; reg_b = prime4; reg_acc = reg_o; o3_X = reg_o; operation : a*b + acc;
"000000100001110000010000100000000000010001110011010111",
--  (425) multiplication_with_reduction_199
-- reg_a = a5_X; reg_b = b6_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001110000000000100000100001000100011010100011",
--  (426) multiplication_with_reduction_200
-- reg_a = o5_X; reg_b = prime6; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100011010110111",
--  (427) multiplication_with_reduction_201
-- reg_a = a6_X; reg_b = b5_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001110000000000100000000000100100010111000011",
--  (428) multiplication_with_reduction_202
-- reg_a = o6_X; reg_b = prime5; reg_acc = reg_o; o4_X = reg_o; operation : a*b + acc;
"000000100001110000010000100000000000010110010111010111",
--  (429) multiplication_with_reduction_203
-- reg_a = a6_X; reg_b = b6_X; reg_acc = reg_o >> 256; Enable sign a, b; operation : a*b + acc;
"000000100001110000000000100000100001100100011011000011",
--  (430) multiplication_with_reduction_204
-- reg_a = o6_X; reg_b = prime6; reg_acc = reg_o; o5_X = reg_o; o6_0 = reg_o >> 256; operation : a*b + acc;
"000000100001110001110000100000000000011010111011010111",
--  (431) multiplication_with_reduction_205
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (432) multiplication_with_reduction_206
-- -- In case of size 8
-- reg_a = a0_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011000000011",
--  (433) multiplication_with_reduction_207
-- reg_a = a6_X; reg_b = b0_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100000011000011",
--  (434) multiplication_with_reduction_208
-- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o6_X = reg_y; operation : keep accumulator;
"000000100001111000011000110000000100011111000000011011",
--  (435) multiplication_with_reduction_209
-- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000010000100000000010011",
--  (436) multiplication_with_reduction_210
-- reg_a = o0_X; reg_b = prime7; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001111000000000100000100000000100011100010111",
--  (437) multiplication_with_reduction_211
-- reg_a = a1_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011000100011",
--  (438) multiplication_with_reduction_212
-- reg_a = o1_X; reg_b = prime6; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011000110111",
--  (439) multiplication_with_reduction_213
-- reg_a = a2_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010101000011",
--  (440) multiplication_with_reduction_214
-- reg_a = o2_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010101010111",
--  (441) multiplication_with_reduction_215
-- reg_a = a3_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010001100011",
--  (442) multiplication_with_reduction_216
-- reg_a = o3_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010001110111",
--  (443) multiplication_with_reduction_217
-- reg_a = a4_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001110000011",
--  (444) multiplication_with_reduction_218
-- reg_a = o4_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001110010111",
--  (445) multiplication_with_reduction_219
-- reg_a = a5_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001010100011",
--  (446) multiplication_with_reduction_220
-- reg_a = o5_X; reg_b = prime2; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001010110111",
--  (447) multiplication_with_reduction_221
-- reg_a = a6_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100000111000011",
--  (448) multiplication_with_reduction_222
-- reg_a = o6_X; reg_b = prime1; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100000111010111",
--  (449) multiplication_with_reduction_223
-- reg_a = a0_X; reg_b = b7_X; reg_acc = reg_o; Enable sign b; operation : a*b + acc;
"000000100001111000000000100000000001000100011100000011",
--  (450) multiplication_with_reduction_224
-- reg_a = a7_X; reg_b = b0_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001111000000000100000000000100100000011100011",
--  (451) multiplication_with_reduction_225
-- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o7_X = reg_y; operation : keep accumulator;
"000000100001111000011000110000000100011111100000011011",
--  (452) multiplication_with_reduction_226
-- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000010000100000000010011",
--  (453) multiplication_with_reduction_227
-- reg_a = a1_X; reg_b = b7_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001111000000000100000100001000100011100100011",
--  (454) multiplication_with_reduction_228
-- reg_a = o1_X; reg_b = prime7; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011100110111",
--  (455) multiplication_with_reduction_229
-- reg_a = a2_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011001000011",
--  (456) multiplication_with_reduction_230
-- reg_a = o2_X; reg_b = prime6; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011001010111",
--  (457) multiplication_with_reduction_231
-- reg_a = a3_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010101100011",
--  (458) multiplication_with_reduction_232
-- reg_a = o3_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010101110111",
--  (459) multiplication_with_reduction_233
-- reg_a = a4_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010010000011",
--  (460) multiplication_with_reduction_234
-- reg_a = o4_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010010010111",
--  (461) multiplication_with_reduction_235
-- reg_a = a5_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001110100011",
--  (462) multiplication_with_reduction_236
-- reg_a = o5_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001110110111",
--  (463) multiplication_with_reduction_237
-- reg_a = a6_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001011000011",
--  (464) multiplication_with_reduction_238
-- reg_a = o6_X; reg_b = prime2; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001011010111",
--  (465) multiplication_with_reduction_239
-- reg_a = a7_X; reg_b = b1_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001111000000000100000000000100100000111100011",
--  (466) multiplication_with_reduction_240
-- reg_a = o7_X; reg_b = prime1; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000000100000111110111",
--  (467) multiplication_with_reduction_241
-- reg_a = a2_X; reg_b = b7_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001111000000000100000100001000100011101000011",
--  (468) multiplication_with_reduction_242
-- reg_a = o2_X; reg_b = prime7; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011101010111",
--  (469) multiplication_with_reduction_243
-- reg_a = a3_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011001100011",
--  (470) multiplication_with_reduction_244
-- reg_a = o3_X; reg_b = prime6; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011001110111",
--  (471) multiplication_with_reduction_245
-- reg_a = a4_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010110000011",
--  (472) multiplication_with_reduction_246
-- reg_a = o4_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010110010111",
--  (473) multiplication_with_reduction_247
-- reg_a = a5_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010010100011",
--  (474) multiplication_with_reduction_248
-- reg_a = o5_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010010110111",
--  (475) multiplication_with_reduction_249
-- reg_a = a6_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001111000011",
--  (476) multiplication_with_reduction_250
-- reg_a = o6_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001111010111",
--  (477) multiplication_with_reduction_251
-- reg_a = a7_X; reg_b = b2_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001111000000000100000000000100100001011100011",
--  (478) multiplication_with_reduction_252
-- reg_a = o7_X; reg_b = prime2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000001000101011110111",
--  (479) multiplication_with_reduction_253
-- reg_a = a3_X; reg_b = b7_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001111000000000100000100001000100011101100011",
--  (480) multiplication_with_reduction_254
-- reg_a = o3_X; reg_b = prime7; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011101110111",
--  (481) multiplication_with_reduction_255
-- reg_a = a4_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011010000011",
--  (482) multiplication_with_reduction_256
-- reg_a = o4_X; reg_b = prime6; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011010010111",
--  (483) multiplication_with_reduction_257
-- reg_a = a5_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010110100011",
--  (484) multiplication_with_reduction_258
-- reg_a = o5_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010110110111",
--  (485) multiplication_with_reduction_259
-- reg_a = a6_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010011000011",
--  (486) multiplication_with_reduction_260
-- reg_a = o6_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010011010111",
--  (487) multiplication_with_reduction_261
-- reg_a = a7_X; reg_b = b3_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001111000000000100000000000100100001111100011",
--  (488) multiplication_with_reduction_262
-- reg_a = o7_X; reg_b = prime3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000001101001111110111",
--  (489) multiplication_with_reduction_263
-- reg_a = a4_X; reg_b = b7_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001111000000000100000100001000100011110000011",
--  (490) multiplication_with_reduction_264
-- reg_a = o4_X; reg_b = prime7; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011110010111",
--  (491) multiplication_with_reduction_265
-- reg_a = a5_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011010100011",
--  (492) multiplication_with_reduction_266
-- reg_a = o5_X; reg_b = prime6; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011010110111",
--  (493) multiplication_with_reduction_267
-- reg_a = a6_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010111000011",
--  (494) multiplication_with_reduction_268
-- reg_a = o6_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010111010111",
--  (495) multiplication_with_reduction_269
-- reg_a = a7_X; reg_b = b4_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001111000000000100000000000100100010011100011",
--  (496) multiplication_with_reduction_270
-- reg_a = o7_X; reg_b = prime4; reg_acc = reg_o; o3_X = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000010001110011110111",
--  (497) multiplication_with_reduction_271
-- reg_a = a5_X; reg_b = b7_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001111000000000100000100001000100011110100011",
--  (498) multiplication_with_reduction_272
-- reg_a = o5_X; reg_b = prime7; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011110110111",
--  (499) multiplication_with_reduction_273
-- reg_a = a6_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011011000011",
--  (500) multiplication_with_reduction_274
-- reg_a = o6_X; reg_b = prime6; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011011010111",
--  (501) multiplication_with_reduction_275
-- reg_a = a7_X; reg_b = b5_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001111000000000100000000000100100010111100011",
--  (502) multiplication_with_reduction_276
-- reg_a = o7_X; reg_b = prime5; reg_acc = reg_o; o4_X = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000010110010111110111",
--  (503) multiplication_with_reduction_277
-- reg_a = a6_X; reg_b = b7_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001111000000000100000100001000100011111000011",
--  (504) multiplication_with_reduction_278
-- reg_a = o6_X; reg_b = prime7; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011111010111",
--  (505) multiplication_with_reduction_279
-- reg_a = a7_X; reg_b = b6_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001111000000000100000000000100100011011100011",
--  (506) multiplication_with_reduction_280
-- reg_a = o7_X; reg_b = prime6; reg_acc = reg_o; o5_X = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000011010111011110111",
--  (507) multiplication_with_reduction_281
-- reg_a = a7_X; reg_b = b7_X; reg_acc = reg_o >> 256; Enable sign a, b; operation : a*b + acc;
"000000100001111000000000100000100001100100011111100011",
--  (508) multiplication_with_reduction_282
-- reg_a = o7_X; reg_b = prime7; reg_acc = reg_o; o6_X = reg_o; o7_0 = reg_o >> 256; operation : a*b + acc;
"000000100001111001110000100000000000011111011111110111",
--  (509) multiplication_with_reduction_283
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (510) multiplication_with_reduction_special_prime_1_0
-- -- In case of size 1
-- reg_a = a0_X; reg_b = b0_X; reg_acc = 0; Enable sign a,b; operation : a*b + acc;
"000000100001000000000000100000010000000100000000000011",
--  (511) multiplication_with_reduction_special_prime_1_1
-- reg_a = 0; reg_b = 0; reg_acc = reg_o >> 256; o0_X = reg_o; operation : a*b + acc;
"000000100001000000010000100000101110000100000000000011",
--  (512) multiplication_with_reduction_special_prime_1_2
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (513) multiplication_with_reduction_special_prime_1_3
-- -- In case of sizes 2, 3, 4, 5, 6, 7, 8
-- reg_a = a0_X; reg_b = b0_X; reg_acc = 0; o0_X = reg_o; operation : a*b + acc;
"000011100001001000010000100000010000000100000000000011",
--  (514) multiplication_with_reduction_special_prime_1_4
-- -- In case of size 2
-- reg_a = a0_X; reg_b = b1_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001001000000000100000100001000100000100000011",
--  (515) multiplication_with_reduction_special_prime_1_5
-- reg_a = o0_X; reg_b = primeSP1; reg_acc = reg_o; operation : a*b + acc;
"000000100001001000000000100000000000000100000100010111",
--  (516) multiplication_with_reduction_special_prime_1_6
-- reg_a = a1_X; reg_b = b0_X; reg_acc = reg_o; o1_X = reg_o; Enable sign a; operation : a*b + acc;
"000000100001001000010000100000000000101000100000100011",
--  (517) multiplication_with_reduction_special_prime_1_7
-- reg_a = a1_X; reg_b = b1_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001001000000000100000100001100100000100100011",
--  (518) multiplication_with_reduction_special_prime_1_8
-- reg_a = o1_X; reg_b = primeSP1; reg_acc = reg_o; o0_X = reg_o; o1_X = reg_o >> 256; operation : a*b + acc;
"000000100001001001110000100000000000000100000100110111",
--  (519) multiplication_with_reduction_special_prime_1_9
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (520) multiplication_with_reduction_special_prime_1_10
-- -- In case of sizes 3, 4, 5, 6, 7, 8
-- reg_a = a0_X; reg_b = b1_X; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001010000000000100000100000000100000100000011",
--  (521) multiplication_with_reduction_special_prime_1_11
-- reg_a = o0_X; reg_b = primeSP1; reg_acc = reg_o; operation : a*b + acc;
"000000100001010000000000100000000000000100000100010111",
--  (522) multiplication_with_reduction_special_prime_1_12
-- reg_a = a1_X; reg_b = b0_X; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
"000000100001010000010000100000000000001000100000100011",
--  (523) multiplication_with_reduction_special_prime_1_13
-- reg_a = o0_X; reg_b = primeSP2; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001010000000000100000100000000100001000010111",
--  (524) multiplication_with_reduction_special_prime_1_14
-- reg_a = a1_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001010000000000100000000000000100000100100011",
--  (525) multiplication_with_reduction_special_prime_1_15
-- reg_a = o1_X; reg_b = primeSP1; reg_acc = reg_o; operation : a*b + acc;
"000101000001010000000000100000000000000100000100110111",
--  (526) multiplication_with_reduction_special_prime_1_16
-- -- In case of size 3
-- reg_a = a0_X; reg_b = b2_X; reg_acc = reg_o; Enable sign b; operation : a*b + acc;
"000000100001010000000000100000000001000100001000000011",
--  (527) multiplication_with_reduction_special_prime_1_17
-- reg_a = a2_X; reg_b = b0_X; reg_acc = reg_o; o2_X = reg_o; Enable sign a; operation : a*b + acc;
"000000100001010000010000100000000000101101000001000011",
--  (528) multiplication_with_reduction_special_prime_1_18
-- reg_a = a1_X; reg_b = b2_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001010000000000100000100001000100001000100011",
--  (529) multiplication_with_reduction_special_prime_1_19
-- reg_a = o1_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
"000000100001010000000000100000000000000100001000110111",
--  (530) multiplication_with_reduction_special_prime_1_20
-- reg_a = a2_X; reg_b = b1_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001010000000000100000000000100100000101000011",
--  (531) multiplication_with_reduction_special_prime_1_21
-- reg_a = o2_X; reg_b = primeSP1; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
"000000100001010000010000100000000000000100000101010111",
--  (532) multiplication_with_reduction_special_prime_1_22
-- reg_a = a2_X; reg_b = b2_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001010000000000100000100001100100001001000011",
--  (533) multiplication_with_reduction_special_prime_1_23
-- reg_a = o2_X; reg_b = primeSP2; reg_acc = reg_o; o1_X = reg_o; o2_X = reg_o >> 256; operation : a*b + acc;
"000000100001010001110000100000000000001000101001010111",
--  (534) multiplication_with_reduction_special_prime_1_24
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (535) multiplication_with_reduction_special_prime_1_25
-- -- In case of sizes 4, 5, 6, 7, 8
-- reg_a = a0_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001011000000000100000000000000100001000000011",
--  (536) multiplication_with_reduction_special_prime_1_26
-- reg_a = a2_X; reg_b = b0_X; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
"000000100001011000010000100000000000001101000001000011",
--  (537) multiplication_with_reduction_special_prime_1_27
-- reg_a = o0_X; reg_b = primeSP3; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001011000000000100000100000000100001100010111",
--  (538) multiplication_with_reduction_special_prime_1_28
-- reg_a = a1_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001011000000000100000000000000100001000100011",
--  (539) multiplication_with_reduction_special_prime_1_29
-- reg_a = o1_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
"000000100001011000000000100000000000000100001000110111",
--  (540) multiplication_with_reduction_special_prime_1_30
-- reg_a = a2_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001011000000000100000000000000100000101000011",
--  (541) multiplication_with_reduction_special_prime_1_31
-- reg_a = o2_X; reg_b = primeSP1; reg_acc = reg_o; operation : a*b + acc;
"001000000001011000000000100000000000000100000101010111",
--  (542) multiplication_with_reduction_special_prime_1_32
-- -- In case of size 4
-- reg_a = a0_X; reg_b = b3_X; reg_acc = reg_o; Enable sign b; operation : a*b + acc;
"000000100001011000000000100000000001000100001100000011",
--  (543) multiplication_with_reduction_special_prime_1_33
-- reg_a = a3_X; reg_b = b0_X; reg_acc = reg_o; o3_X = reg_o; Enable sign a; operation : a*b + acc;
"000000100001011000010000100000000000100001100001100011",
--  (544) multiplication_with_reduction_special_prime_1_34
-- reg_a = a1_X; reg_b = b3_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001011000000000100000100001000100001100100011",
--  (545) multiplication_with_reduction_special_prime_1_35
-- reg_a = o1_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001011000000000100000000000000100001100110111",
--  (546) multiplication_with_reduction_special_prime_1_36
-- reg_a = a2_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001011000000000100000000000000100001001000011",
--  (547) multiplication_with_reduction_special_prime_1_37
-- reg_a = o2_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
"000000100001011000000000100000000000000100001001010111",
--  (548) multiplication_with_reduction_special_prime_1_38
-- reg_a = a3_X; reg_b = b1_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001011000000000100000000000100100000101100011",
--  (549) multiplication_with_reduction_special_prime_1_39
-- reg_a = o3_X; reg_b = primeSP1; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
"000000100001011000010000100000000000000100000101110111",
--  (550) multiplication_with_reduction_special_prime_1_40
-- reg_a = a2_X; reg_b = b3_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001011000000000100000100001000100001101000011",
--  (551) multiplication_with_reduction_special_prime_1_41
-- reg_a = o2_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001011000000000100000000000000100001101010111",
--  (552) multiplication_with_reduction_special_prime_1_42
-- reg_a = a3_X; reg_b = b2_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001011000000000100000000000100100001001100011",
--  (553) multiplication_with_reduction_special_prime_1_43
-- reg_a = o3_X; reg_b = primeSP2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
"000000100001011000010000100000000000001000101001110111",
--  (554) multiplication_with_reduction_special_prime_1_44
-- reg_a = a3_X; reg_b = b3_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001011000000000100000100001100100001101100011",
--  (555) multiplication_with_reduction_special_prime_1_45
-- reg_a = o3_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; o3_X = reg_o >> 256; operation : a*b + acc;
"000000100001011001110000100000000000001101001101110111",
--  (556) multiplication_with_reduction_special_prime_1_46
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (557) multiplication_with_reduction_special_prime_1_47
-- -- In case of sizes 5, 6, 7, 8
-- reg_a = a0_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001100000011",
--  (558) multiplication_with_reduction_special_prime_1_48
-- reg_a = a3_X; reg_b = b0_X; reg_acc = reg_o; o3_X = reg_o; operation : a*b + acc;
"000000100001100000010000100000000000010001100001100011",
--  (559) multiplication_with_reduction_special_prime_1_49
-- reg_a = o0_X; reg_b = primeSP4; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001100000000000100000100000000100010000010111",
--  (560) multiplication_with_reduction_special_prime_1_50
-- reg_a = a1_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001100100011",
--  (561) multiplication_with_reduction_special_prime_1_51
-- reg_a = o1_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001100110111",
--  (562) multiplication_with_reduction_special_prime_1_52
-- reg_a = a2_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001001000011",
--  (563) multiplication_with_reduction_special_prime_1_53
-- reg_a = o2_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001001010111",
--  (564) multiplication_with_reduction_special_prime_1_54
-- reg_a = a3_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100000101100011",
--  (565) multiplication_with_reduction_special_prime_1_55
-- reg_a = o3_X; reg_b = primeSP1; reg_acc = reg_o; operation : a*b + acc;
"001100000001100000000000100000000000000100000101110111",
--  (566) multiplication_with_reduction_special_prime_1_56
-- -- In case of size 5
-- reg_a = a0_X; reg_b = b4_X; reg_acc = reg_o; Enable sign b; operation : a*b + acc;
"000000100001100000000000100000000001000100010000000011",
--  (567) multiplication_with_reduction_special_prime_1_57
-- reg_a = a4_X; reg_b = b0_X; reg_acc = reg_o; o4_X = reg_o; Enable sign a; operation : a*b + acc;
"000000100001100000010000100000000000110110000010000011",
--  (568) multiplication_with_reduction_special_prime_1_58
-- reg_a = a1_X; reg_b = b4_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001100000000000100000100001000100010000100011",
--  (569) multiplication_with_reduction_special_prime_1_59
-- reg_a = o1_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100010000110111",
--  (570) multiplication_with_reduction_special_prime_1_60
-- reg_a = a2_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001101000011",
--  (571) multiplication_with_reduction_special_prime_1_61
-- reg_a = o2_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001101010111",
--  (572) multiplication_with_reduction_special_prime_1_62
-- reg_a = a3_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001001100011",
--  (573) multiplication_with_reduction_special_prime_1_63
-- reg_a = o3_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001001110111",
--  (574) multiplication_with_reduction_special_prime_1_64
-- reg_a = a4_X; reg_b = b1_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001100000000000100000000000100100000110000011",
--  (575) multiplication_with_reduction_special_prime_1_65
-- reg_a = o4_X; reg_b = primeSP1; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
"000000100001100000010000100000000000000100000110010111",
--  (576) multiplication_with_reduction_special_prime_1_66
-- reg_a = a2_X; reg_b = b4_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001100000000000100000100001000100010001000011",
--  (577) multiplication_with_reduction_special_prime_1_67
-- reg_a = o2_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100010001010111",
--  (578) multiplication_with_reduction_special_prime_1_68
-- reg_a = a3_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001101100011",
--  (579) multiplication_with_reduction_special_prime_1_69
-- reg_a = o3_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001101110111",
--  (580) multiplication_with_reduction_special_prime_1_70
-- reg_a = a4_X; reg_b = b2_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001100000000000100000000000100100001010000011",
--  (581) multiplication_with_reduction_special_prime_1_71
-- reg_a = o4_X; reg_b = primeSP2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
"000000100001100000010000100000000000001000101010010111",
--  (582) multiplication_with_reduction_special_prime_1_72
-- reg_a = a3_X; reg_b = b4_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001100000000000100000100001000100010001100011",
--  (583) multiplication_with_reduction_special_prime_1_73
-- reg_a = o3_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100010001110111",
--  (584) multiplication_with_reduction_special_prime_1_74
-- reg_a = a4_X; reg_b = b3_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001100000000000100000000000100100001110000011",
--  (585) multiplication_with_reduction_special_prime_1_75
-- reg_a = o4_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
"000000100001100000010000100000000000001101001110010111",
--  (586) multiplication_with_reduction_special_prime_1_76
-- reg_a = a4_X; reg_b = b4_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001100000000000100000100001100100010010000011",
--  (587) multiplication_with_reduction_special_prime_1_77
-- reg_a = o4_X; reg_b = primeSP4; reg_acc = reg_o; o3_X = reg_o; o4_X = reg_o >> 256; operation : a*b + acc;
"000000100001100001110000100000000000010001110010010111",
--  (588) multiplication_with_reduction_special_prime_1_78
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (589) multiplication_with_reduction_special_prime_1_79
-- -- In case of sizes 6, 7, 8
-- reg_a = a0_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010000000011",
--  (590) multiplication_with_reduction_special_prime_1_80
-- reg_a = a4_X; reg_b = b0_X; reg_acc = reg_o; o4_X = reg_o; operation : a*b + acc;
"000000100001101000010000100000000000010110000010000011",
--  (591) multiplication_with_reduction_special_prime_1_81
-- reg_a = o0_X; reg_b = primeSP5; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001101000000000100000100000000100010100010111",
--  (592) multiplication_with_reduction_special_prime_1_82
-- reg_a = a1_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010000100011",
--  (593) multiplication_with_reduction_special_prime_1_83
-- reg_a = o1_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010000110111",
--  (594) multiplication_with_reduction_special_prime_1_84
-- reg_a = a2_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001101000011",
--  (595) multiplication_with_reduction_special_prime_1_85
-- reg_a = o2_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001101010111",
--  (596) multiplication_with_reduction_special_prime_1_86
-- reg_a = a3_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001001100011",
--  (597) multiplication_with_reduction_special_prime_1_87
-- reg_a = o3_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001001110111",
--  (598) multiplication_with_reduction_special_prime_1_88
-- reg_a = a4_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100000110000011",
--  (599) multiplication_with_reduction_special_prime_1_89
-- reg_a = o4_X; reg_b = primeSP1; reg_acc = reg_o; operation : a*b + acc;
"010001000001101000000000100000000000000100000110010111",
--  (600) multiplication_with_reduction_special_prime_1_90
-- -- In case of size 6
-- reg_a = a0_X; reg_b = b5_X; reg_acc = reg_o; Enable sign b; operation : a*b + acc;
"000000100001101000000000100000000001000100010100000011",
--  (601) multiplication_with_reduction_special_prime_1_91
-- reg_a = a5_X; reg_b = b0_X; reg_acc = reg_o; o5_X = reg_o; Enable sign a; operation : a*b + acc;
"000000100001101000010000100000000000111010100010100011",
--  (602) multiplication_with_reduction_special_prime_1_92
-- reg_a = a1_X; reg_b = b5_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001101000000000100000100001000100010100100011",
--  (603) multiplication_with_reduction_special_prime_1_93
-- reg_a = o1_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010100110111",
--  (604) multiplication_with_reduction_special_prime_1_94
-- reg_a = a2_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010001000011",
--  (605) multiplication_with_reduction_special_prime_1_95
-- reg_a = o2_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010001010111",
--  (606) multiplication_with_reduction_special_prime_1_96
-- reg_a = a3_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001101100011",
--  (607) multiplication_with_reduction_special_prime_1_97
-- reg_a = o3_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001101110111",
--  (608) multiplication_with_reduction_special_prime_1_98
-- reg_a = a4_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001010000011",
--  (609) multiplication_with_reduction_special_prime_1_99
-- reg_a = o4_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001010010111",
--  (610) multiplication_with_reduction_special_prime_1_100
-- reg_a = a5_X; reg_b = b1_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001101000000000100000000000100100000110100011",
--  (611) multiplication_with_reduction_special_prime_1_101
-- reg_a = o5_X; reg_b = primeSP1; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
"000000100001101000010000100000000000000100000110110111",
--  (612) multiplication_with_reduction_special_prime_1_102
-- reg_a = a2_X; reg_b = b5_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001101000000000100000100001000100010101000011",
--  (613) multiplication_with_reduction_special_prime_1_103
-- reg_a = o2_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010101010111",
--  (614) multiplication_with_reduction_special_prime_1_104
-- reg_a = a3_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010001100011",
--  (615) multiplication_with_reduction_special_prime_1_105
-- reg_a = o3_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010001110111",
--  (616) multiplication_with_reduction_special_prime_1_106
-- reg_a = a4_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001110000011",
--  (617) multiplication_with_reduction_special_prime_1_107
-- reg_a = o4_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001110010111",
--  (618) multiplication_with_reduction_special_prime_1_108
-- reg_a = a5_X; reg_b = b2_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001101000000000100000000000100100001010100011",
--  (619) multiplication_with_reduction_special_prime_1_109
-- reg_a = o5_X; reg_b = primeSP2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
"000000100001101000010000100000000000001000101010110111",
--  (620) multiplication_with_reduction_special_prime_1_110
-- reg_a = a3_X; reg_b = b5_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001101000000000100000100001000100010101100011",
--  (621) multiplication_with_reduction_special_prime_1_111
-- reg_a = o3_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010101110111",
--  (622) multiplication_with_reduction_special_prime_1_112
-- reg_a = a4_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010010000011",
--  (623) multiplication_with_reduction_special_prime_1_113
-- reg_a = o4_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010010010111",
--  (624) multiplication_with_reduction_special_prime_1_114
-- reg_a = a5_X; reg_b = b3_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001101000000000100000000000100100001110100011",
--  (625) multiplication_with_reduction_special_prime_1_115
-- reg_a = o5_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
"000000100001101000010000100000000000001101001110110111",
--  (626) multiplication_with_reduction_special_prime_1_116
-- reg_a = a4_X; reg_b = b5_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001101000000000100000100001000100010110000011",
--  (627) multiplication_with_reduction_special_prime_1_117
-- reg_a = o4_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010110010111",
--  (628) multiplication_with_reduction_special_prime_1_118
-- reg_a = a5_X; reg_b = b4_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001101000000000100000000000100100010010100011",
--  (629) multiplication_with_reduction_special_prime_1_119
-- reg_a = o5_X; reg_b = primeSP4; reg_acc = reg_o; o3_X = reg_o; operation : a*b + acc;
"000000100001101000010000100000000000010001110010110111",
--  (630) multiplication_with_reduction_special_prime_1_120
-- reg_a = a5_X; reg_b = b5_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001101000000000100000100001100100010110100011",
--  (631) multiplication_with_reduction_special_prime_1_121
-- reg_a = o5_X; reg_b = primeSP5; reg_acc = reg_o; o4_X = reg_o; o5_X = reg_o >> 256; operation : a*b + acc;
"000000100001101001110000100000000000010110010110110111",
--  (632) multiplication_with_reduction_special_prime_1_122
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (633) multiplication_with_reduction_special_prime_1_123
-- -- In case of sizes 7, 8
-- reg_a = a0_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010100000011",
--  (634) multiplication_with_reduction_special_prime_1_124
-- reg_a = a5_X; reg_b = b0_X; reg_acc = reg_o; o5_X = reg_o; operation : a*b + acc;
"000000100001110000010000100000000000011010100010100011",
--  (635) multiplication_with_reduction_special_prime_1_125
-- reg_a = o0_X; reg_b = primeSP6; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001110000000000100000100000000100011000010111",
--  (636) multiplication_with_reduction_special_prime_1_126
-- reg_a = a1_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010100100011",
--  (637) multiplication_with_reduction_special_prime_1_127
-- reg_a = o1_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010100110111",
--  (638) multiplication_with_reduction_special_prime_1_128
-- reg_a = a2_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010001000011",
--  (639) multiplication_with_reduction_special_prime_1_129
-- reg_a = o2_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010001010111",
--  (640) multiplication_with_reduction_special_prime_1_130
-- reg_a = a3_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001101100011",
--  (641) multiplication_with_reduction_special_prime_1_131
-- reg_a = o3_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001101110111",
--  (642) multiplication_with_reduction_special_prime_1_132
-- reg_a = a4_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001010000011",
--  (643) multiplication_with_reduction_special_prime_1_133
-- reg_a = o4_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001010010111",
--  (644) multiplication_with_reduction_special_prime_1_134
-- reg_a = a5_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100000110100011",
--  (645) multiplication_with_reduction_special_prime_1_135
-- reg_a = o5_X; reg_b = primeSP1; reg_acc = reg_o; operation : a*b + acc;
"010111000001110000000000100000000000000100000110110111",
--  (646) multiplication_with_reduction_special_prime_1_136
-- -- In case of size 7
-- reg_a = a0_X; reg_b = b6_X; reg_acc = reg_o; Enable sign b; operation : a*b + acc;
"000000100001110000000000100000000001000100011000000011",
--  (647) multiplication_with_reduction_special_prime_1_137
-- reg_a = a6_X; reg_b = b0_X; reg_acc = reg_o; o6_X = reg_o; Enable sign a; operation : a*b + acc;
"000000100001110000010000100000000000111111000011000011",
--  (648) multiplication_with_reduction_special_prime_1_138
-- reg_a = a1_X; reg_b = b6_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001110000000000100000100001000100011000100011",
--  (649) multiplication_with_reduction_special_prime_1_139
-- reg_a = o1_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100011000110111",
--  (650) multiplication_with_reduction_special_prime_1_140
-- reg_a = a2_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010101000011",
--  (651) multiplication_with_reduction_special_prime_1_141
-- reg_a = o2_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010101010111",
--  (652) multiplication_with_reduction_special_prime_1_142
-- reg_a = a3_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010001100011",
--  (653) multiplication_with_reduction_special_prime_1_143
-- reg_a = o3_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010001110111",
--  (654) multiplication_with_reduction_special_prime_1_144
-- reg_a = a4_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001110000011",
--  (655) multiplication_with_reduction_special_prime_1_145
-- reg_a = o4_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001110010111",
--  (656) multiplication_with_reduction_special_prime_1_146
-- reg_a = a5_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001010100011",
--  (657) multiplication_with_reduction_special_prime_1_147
-- reg_a = o5_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001010110111",
--  (658) multiplication_with_reduction_special_prime_1_148
-- reg_a = a6_X; reg_b = b1_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001110000000000100000000000100100000111000011",
--  (659) multiplication_with_reduction_special_prime_1_149
-- reg_a = o6_X; reg_b = primeSP1; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
"000000100001110000010000100000000000000100000111010111",
--  (660) multiplication_with_reduction_special_prime_1_150
-- reg_a = a2_X; reg_b = b6_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001110000000000100000100001000100011001000011",
--  (661) multiplication_with_reduction_special_prime_1_151
-- reg_a = o2_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100011001010111",
--  (662) multiplication_with_reduction_special_prime_1_152
-- reg_a = a3_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010101100011",
--  (663) multiplication_with_reduction_special_prime_1_153
-- reg_a = o3_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010101110111",
--  (664) multiplication_with_reduction_special_prime_1_154
-- reg_a = a4_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010010000011",
--  (665) multiplication_with_reduction_special_prime_1_155
-- reg_a = o4_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010010010111",
--  (666) multiplication_with_reduction_special_prime_1_156
-- reg_a = a5_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001110100011",
--  (667) multiplication_with_reduction_special_prime_1_157
-- reg_a = o5_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001110110111",
--  (668) multiplication_with_reduction_special_prime_1_158
-- reg_a = a6_X; reg_b = b2_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001110000000000100000000000100100001011000011",
--  (669) multiplication_with_reduction_special_prime_1_159
-- reg_a = o6_X; reg_b = primeSP2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
"000000100001110000010000100000000000001000101011010111",
--  (670) multiplication_with_reduction_special_prime_1_160
-- reg_a = a3_X; reg_b = b6_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001110000000000100000100001000100011001100011",
--  (671) multiplication_with_reduction_special_prime_1_161
-- reg_a = o3_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100011001110111",
--  (672) multiplication_with_reduction_special_prime_1_162
-- reg_a = a4_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010110000011",
--  (673) multiplication_with_reduction_special_prime_1_163
-- reg_a = o4_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010110010111",
--  (674) multiplication_with_reduction_special_prime_1_164
-- reg_a = a5_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010010100011",
--  (675) multiplication_with_reduction_special_prime_1_165
-- reg_a = o5_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010010110111",
--  (676) multiplication_with_reduction_special_prime_1_166
-- reg_a = a6_X; reg_b = b3_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001110000000000100000000000100100001111000011",
--  (677) multiplication_with_reduction_special_prime_1_167
-- reg_a = o6_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
"000000100001110000010000100000000000001101001111010111",
--  (678) multiplication_with_reduction_special_prime_1_168
-- reg_a = a4_X; reg_b = b6_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001110000000000100000100001000100011010000011",
--  (679) multiplication_with_reduction_special_prime_1_169
-- reg_a = o4_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100011010010111",
--  (680) multiplication_with_reduction_special_prime_1_170
-- reg_a = a5_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010110100011",
--  (681) multiplication_with_reduction_special_prime_1_171
-- reg_a = o5_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010110110111",
--  (682) multiplication_with_reduction_special_prime_1_172
-- reg_a = a6_X; reg_b = b4_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001110000000000100000000000100100010011000011",
--  (683) multiplication_with_reduction_special_prime_1_173
-- reg_a = o6_X; reg_b = primeSP4; reg_acc = reg_o; o3_X = reg_o; operation : a*b + acc;
"000000100001110000010000100000000000010001110011010111",
--  (684) multiplication_with_reduction_special_prime_1_174
-- reg_a = a5_X; reg_b = b6_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001110000000000100000100001000100011010100011",
--  (685) multiplication_with_reduction_special_prime_1_175
-- reg_a = o5_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100011010110111",
--  (686) multiplication_with_reduction_special_prime_1_176
-- reg_a = a6_X; reg_b = b5_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001110000000000100000000000100100010111000011",
--  (687) multiplication_with_reduction_special_prime_1_177
-- reg_a = o6_X; reg_b = primeSP5; reg_acc = reg_o; o4_X = reg_o; operation : a*b + acc;
"000000100001110000010000100000000000010110010111010111",
--  (688) multiplication_with_reduction_special_prime_1_178
-- reg_a = a6_X; reg_b = b6_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001110000000000100000100001100100011011000011",
--  (689) multiplication_with_reduction_special_prime_1_179
-- reg_a = o6_X; reg_b = primeSP6; reg_acc = reg_o; o5_X = reg_o; o6_X = reg_o >> 256; operation : a*b + acc;
"000000100001110001110000100000000000011010111011010111",
--  (690) multiplication_with_reduction_special_prime_1_180
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (691) multiplication_with_reduction_special_prime_1_181
-- -- In case of size 8
-- reg_a = a0_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011000000011",
--  (692) multiplication_with_reduction_special_prime_1_182
-- reg_a = a6_X; reg_b = b0_X; reg_acc = reg_o; o6_X = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000011111000011000011",
--  (693) multiplication_with_reduction_special_prime_1_183
-- reg_a = o0_X; reg_b = primeSP7; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001111000000000100000100000000100011100010111",
--  (694) multiplication_with_reduction_special_prime_1_184
-- reg_a = a1_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011000100011",
--  (695) multiplication_with_reduction_special_prime_1_185
-- reg_a = o1_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011000110111",
--  (696) multiplication_with_reduction_special_prime_1_186
-- reg_a = a2_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010101000011",
--  (697) multiplication_with_reduction_special_prime_1_187
-- reg_a = o2_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010101010111",
--  (698) multiplication_with_reduction_special_prime_1_188
-- reg_a = a3_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010001100011",
--  (699) multiplication_with_reduction_special_prime_1_189
-- reg_a = o3_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010001110111",
--  (700) multiplication_with_reduction_special_prime_1_190
-- reg_a = a4_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001110000011",
--  (701) multiplication_with_reduction_special_prime_1_191
-- reg_a = o4_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001110010111",
--  (702) multiplication_with_reduction_special_prime_1_192
-- reg_a = a5_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001010100011",
--  (703) multiplication_with_reduction_special_prime_1_193
-- reg_a = o5_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001010110111",
--  (704) multiplication_with_reduction_special_prime_1_194
-- reg_a = a6_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100000111000011",
--  (705) multiplication_with_reduction_special_prime_1_195
-- reg_a = o6_X; reg_b = primeSP1; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100000111010111",
--  (706) multiplication_with_reduction_special_prime_1_196
-- reg_a = a0_X; reg_b = b7_X; reg_acc = reg_o; Enable sign b; operation : a*b + acc;
"000000100001111000000000100000000001000100011100000011",
--  (707) multiplication_with_reduction_special_prime_1_197
-- reg_a = a7_X; reg_b = b0_X; reg_acc = reg_o; o7_X = reg_o; Enable sign a; operation : a*b + acc;
"000000100001111000010000100000000000100011100011100011",
--  (708) multiplication_with_reduction_special_prime_1_198
-- reg_a = a1_X; reg_b = b7_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001111000000000100000100001000100011100100011",
--  (709) multiplication_with_reduction_special_prime_1_199
-- reg_a = o1_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011100110111",
--  (710) multiplication_with_reduction_special_prime_1_200
-- reg_a = a2_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011001000011",
--  (711) multiplication_with_reduction_special_prime_1_201
-- reg_a = o2_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011001010111",
--  (712) multiplication_with_reduction_special_prime_1_202
-- reg_a = a3_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010101100011",
--  (713) multiplication_with_reduction_special_prime_1_203
-- reg_a = o3_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010101110111",
--  (714) multiplication_with_reduction_special_prime_1_204
-- reg_a = a4_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010010000011",
--  (715) multiplication_with_reduction_special_prime_1_205
-- reg_a = o4_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010010010111",
--  (716) multiplication_with_reduction_special_prime_1_206
-- reg_a = a5_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001110100011",
--  (717) multiplication_with_reduction_special_prime_1_207
-- reg_a = o5_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001110110111",
--  (718) multiplication_with_reduction_special_prime_1_208
-- reg_a = a6_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001011000011",
--  (719) multiplication_with_reduction_special_prime_1_209
-- reg_a = o6_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001011010111",
--  (720) multiplication_with_reduction_special_prime_1_210
-- reg_a = a7_X; reg_b = b1_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001111000000000100000000000100100000111100011",
--  (721) multiplication_with_reduction_special_prime_1_211
-- reg_a = o7_X; reg_b = primeSP1; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000000100000111110111",
--  (722) multiplication_with_reduction_special_prime_1_212
-- reg_a = a2_X; reg_b = b7_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001111000000000100000100001000100011101000011",
--  (723) multiplication_with_reduction_special_prime_1_213
-- reg_a = o2_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011101010111",
--  (724) multiplication_with_reduction_special_prime_1_214
-- reg_a = a3_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011001100011",
--  (725) multiplication_with_reduction_special_prime_1_215
-- reg_a = o3_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011001110111",
--  (726) multiplication_with_reduction_special_prime_1_216
-- reg_a = a4_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010110000011",
--  (727) multiplication_with_reduction_special_prime_1_217
-- reg_a = o4_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010110010111",
--  (728) multiplication_with_reduction_special_prime_1_218
-- reg_a = a5_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010010100011",
--  (729) multiplication_with_reduction_special_prime_1_219
-- reg_a = o5_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010010110111",
--  (730) multiplication_with_reduction_special_prime_1_220
-- reg_a = a6_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001111000011",
--  (731) multiplication_with_reduction_special_prime_1_221
-- reg_a = o6_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001111010111",
--  (732) multiplication_with_reduction_special_prime_1_222
-- reg_a = a7_X; reg_b = b2_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001111000000000100000000000100100001011100011",
--  (733) multiplication_with_reduction_special_prime_1_223
-- reg_a = o7_X; reg_b = primeSP2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000001000101011110111",
--  (734) multiplication_with_reduction_special_prime_1_224
-- reg_a = a3_X; reg_b = b7_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001111000000000100000100001000100011101100011",
--  (735) multiplication_with_reduction_special_prime_1_225
-- reg_a = o3_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011101110111",
--  (736) multiplication_with_reduction_special_prime_1_226
-- reg_a = a4_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011010000011",
--  (737) multiplication_with_reduction_special_prime_1_227
-- reg_a = o4_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011010010111",
--  (738) multiplication_with_reduction_special_prime_1_228
-- reg_a = a5_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010110100011",
--  (739) multiplication_with_reduction_special_prime_1_229
-- reg_a = o5_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010110110111",
--  (740) multiplication_with_reduction_special_prime_1_230
-- reg_a = a6_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010011000011",
--  (741) multiplication_with_reduction_special_prime_1_231
-- reg_a = o6_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010011010111",
--  (742) multiplication_with_reduction_special_prime_1_232
-- reg_a = a7_X; reg_b = b3_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001111000000000100000000000100100001111100011",
--  (743) multiplication_with_reduction_special_prime_1_233
-- reg_a = o7_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000001101001111110111",
--  (744) multiplication_with_reduction_special_prime_1_234
-- reg_a = a4_X; reg_b = b7_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001111000000000100000100001000100011110000011",
--  (745) multiplication_with_reduction_special_prime_1_235
-- reg_a = o4_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011110010111",
--  (746) multiplication_with_reduction_special_prime_1_236
-- reg_a = a5_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011010100011",
--  (747) multiplication_with_reduction_special_prime_1_237
-- reg_a = o5_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011010110111",
--  (748) multiplication_with_reduction_special_prime_1_238
-- reg_a = a6_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010111000011",
--  (749) multiplication_with_reduction_special_prime_1_239
-- reg_a = o6_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010111010111",
--  (750) multiplication_with_reduction_special_prime_1_240
-- reg_a = a7_X; reg_b = b4_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001111000000000100000000000100100010011100011",
--  (751) multiplication_with_reduction_special_prime_1_241
-- reg_a = o7_X; reg_b = primeSP4; reg_acc = reg_o; o3_X = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000010001110011110111",
--  (752) multiplication_with_reduction_special_prime_1_242
-- reg_a = a5_X; reg_b = b7_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001111000000000100000100001000100011110100011",
--  (753) multiplication_with_reduction_special_prime_1_243
-- reg_a = o5_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011110110111",
--  (754) multiplication_with_reduction_special_prime_1_244
-- reg_a = a6_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011011000011",
--  (755) multiplication_with_reduction_special_prime_1_245
-- reg_a = o6_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011011010111",
--  (756) multiplication_with_reduction_special_prime_1_246
-- reg_a = a7_X; reg_b = b5_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001111000000000100000000000100100010111100011",
--  (757) multiplication_with_reduction_special_prime_1_247
-- reg_a = o7_X; reg_b = primeSP5; reg_acc = reg_o; o4_X = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000010110010111110111",
--  (758) multiplication_with_reduction_special_prime_1_248
-- reg_a = a6_X; reg_b = b7_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001111000000000100000100001000100011111000011",
--  (759) multiplication_with_reduction_special_prime_1_249
-- reg_a = o6_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011111010111",
--  (760) multiplication_with_reduction_special_prime_1_250
-- reg_a = a7_X; reg_b = b6_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001111000000000100000000000100100011011100011",
--  (761) multiplication_with_reduction_special_prime_1_251
-- reg_a = o7_X; reg_b = primeSP6; reg_acc = reg_o; o5_X = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000011010111011110111",
--  (762) multiplication_with_reduction_special_prime_1_252
-- reg_a = a7_X; reg_b = b7_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001111000000000100000100001100100011111100011",
--  (763) multiplication_with_reduction_special_prime_1_253
-- reg_a = o7_X; reg_b = primeSP7; reg_acc = reg_o; o6_X = reg_o; o7_X = reg_o >> 256; operation : a*b + acc;
"000000100001111001110000100000000000011111011111110111",
--  (764) multiplication_with_reduction_special_prime_1_254
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (765) multiplication_with_reduction_special_prime_2_0
-- With 2 zeroes in prime sharp
-- -- In case of sizes 2, 3, 4, 5, 6, 7, 8
-- reg_a = a0_X; reg_b = b0_X; reg_acc = 0; o0_X = reg_o; operation : a*b + acc;
"000010100001001000010000100000010000000100000000000011",
--  (766) multiplication_with_reduction_special_prime_2_1
-- -- In case of size 2
-- reg_a = a0_X; reg_b = b1_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001001000000000100000100001000100000100000011",
--  (767) multiplication_with_reduction_special_prime_2_2
-- reg_a = a1_X; reg_b = b0_X; reg_acc = reg_o; o1_X = reg_o; Enable sign a; operation : a*b + acc;
"000000100001001000010000100000000000101000100000100011",
--  (768) multiplication_with_reduction_special_prime_2_3
-- reg_a = a1_X; reg_b = b1_X; reg_acc = reg_o >> 256; o0_X = reg_o; o1_X = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001001001110000100000100001100100000100100011",
--  (769) multiplication_with_reduction_special_prime_2_4
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (770) multiplication_with_reduction_special_prime_2_5
-- -- In case of sizes 3, 4, 5, 6, 7, 8
-- reg_a = a0_X; reg_b = b1_X; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001010000000000100000100000000100000100000011",
--  (771) multiplication_with_reduction_special_prime_2_6
-- reg_a = a1_X; reg_b = b0_X; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
"000000100001010000010000100000000000001000100000100011",
--  (772) multiplication_with_reduction_special_prime_2_7
-- reg_a = o0_X; reg_b = primeSP2; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001010000000000100000100000000100001000010111",
--  (773) multiplication_with_reduction_special_prime_2_8
-- reg_a = a1_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
"000100100001010000000000100000000000000100000100100011",
--  (774) multiplication_with_reduction_special_prime_2_9
-- -- In case of size 3
-- reg_a = a0_X; reg_b = b2_X; reg_acc = reg_o; Enable sign b; operation : a*b + acc;
"000000100001010000000000100000000001000100001000000011",
--  (775) multiplication_with_reduction_special_prime_2_10
-- reg_a = a2_X; reg_b = b0_X; reg_acc = reg_o; o2_X = reg_o; Enable sign a; operation : a*b + acc;
"000000100001010000010000100000000000101101000001000011",
--  (776) multiplication_with_reduction_special_prime_2_11
-- reg_a = a1_X; reg_b = b2_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001010000000000100000100001000100001000100011",
--  (777) multiplication_with_reduction_special_prime_2_12
-- reg_a = o1_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
"000000100001010000000000100000000000000100001000110111",
--  (778) multiplication_with_reduction_special_prime_2_13
-- reg_a = a2_X; reg_b = b1_X; reg_acc = reg_o; Enable sign a; o0_X = reg_o; operation : a*b + acc;
"000000100001010000010000100000000000100100000101000011",
--  (779) multiplication_with_reduction_special_prime_2_14
-- reg_a = a2_X; reg_b = b2_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001010000000000100000100001100100001001000011",
--  (780) multiplication_with_reduction_special_prime_2_15
-- reg_a = o2_X; reg_b = primeSP2; reg_acc = reg_o; o1_X = reg_o; o2_X = reg_o >> 256; operation : a*b + acc;
"000000100001010001110000100000000000001000101001010111",
--  (781) multiplication_with_reduction_special_prime_2_16
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (782) multiplication_with_reduction_special_prime_2_17
-- -- In case of sizes 4, 5, 6, 7, 8
-- reg_a = a0_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001011000000000100000000000000100001000000011",
--  (783) multiplication_with_reduction_special_prime_2_18
-- reg_a = a2_X; reg_b = b0_X; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
"000000100001011000010000100000000000001101000001000011",
--  (784) multiplication_with_reduction_special_prime_2_19
-- reg_a = o0_X; reg_b = primeSP3; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001011000000000100000100000000100001100010111",
--  (785) multiplication_with_reduction_special_prime_2_20
-- reg_a = a1_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001011000000000100000000000000100001000100011",
--  (786) multiplication_with_reduction_special_prime_2_21
-- reg_a = o1_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
"000000100001011000000000100000000000000100001000110111",
--  (787) multiplication_with_reduction_special_prime_2_22
-- reg_a = a2_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
"000111100001011000000000100000000000000100000101000011",
--  (788) multiplication_with_reduction_special_prime_2_23
-- -- In case of size 4
-- reg_a = a0_X; reg_b = b3_X; reg_acc = reg_o; Enable sign b; operation : a*b + acc;
"000000100001011000000000100000000001000100001100000011",
--  (789) multiplication_with_reduction_special_prime_2_24
-- reg_a = a3_X; reg_b = b0_X; reg_acc = reg_o; o3_X = reg_o; Enable sign a; operation : a*b + acc;
"000000100001011000010000100000000000100001100001100011",
--  (790) multiplication_with_reduction_special_prime_2_25
-- reg_a = a1_X; reg_b = b3_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001011000000000100000100001000100001100100011",
--  (791) multiplication_with_reduction_special_prime_2_26
-- reg_a = o1_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001011000000000100000000000000100001100110111",
--  (792) multiplication_with_reduction_special_prime_2_27
-- reg_a = a2_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001011000000000100000000000000100001001000011",
--  (793) multiplication_with_reduction_special_prime_2_28
-- reg_a = o2_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
"000000100001011000000000100000000000000100001001010111",
--  (794) multiplication_with_reduction_special_prime_2_29
-- reg_a = a3_X; reg_b = b1_X; reg_acc = reg_o; Enable sign a; o0_X = reg_o; operation : a*b + acc;
"000000100001011000010000100000000000100100000101100011",
--  (795) multiplication_with_reduction_special_prime_2_30
-- reg_a = a2_X; reg_b = b3_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001011000000000100000100001000100001101000011",
--  (796) multiplication_with_reduction_special_prime_2_31
-- reg_a = o2_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001011000000000100000000000000100001101010111",
--  (797) multiplication_with_reduction_special_prime_2_32
-- reg_a = a3_X; reg_b = b2_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001011000000000100000000000100100001001100011",
--  (798) multiplication_with_reduction_special_prime_2_33
-- reg_a = o3_X; reg_b = primeSP2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
"000000100001011000010000100000000000001000101001110111",
--  (799) multiplication_with_reduction_special_prime_2_34
-- reg_a = a3_X; reg_b = b3_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001011000000000100000100001100100001101100011",
--  (800) multiplication_with_reduction_special_prime_2_35
-- reg_a = o3_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; o3_X = reg_o >> 256; operation : a*b + acc;
"000000100001011001110000100000000000001101001101110111",
--  (801) multiplication_with_reduction_special_prime_2_36
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (802) multiplication_with_reduction_special_prime_2_37
-- -- In case of sizes 5, 6, 7, 8
-- reg_a = a0_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001100000011",
--  (803) multiplication_with_reduction_special_prime_2_38
-- reg_a = a3_X; reg_b = b0_X; reg_acc = reg_o; o3_X = reg_o; operation : a*b + acc;
"000000100001100000010000100000000000010001100001100011",
--  (804) multiplication_with_reduction_special_prime_2_39
-- reg_a = o0_X; reg_b = primeSP4; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001100000000000100000100000000100010000010111",
--  (805) multiplication_with_reduction_special_prime_2_40
-- reg_a = a1_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001100100011",
--  (806) multiplication_with_reduction_special_prime_2_41
-- reg_a = o1_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001100110111",
--  (807) multiplication_with_reduction_special_prime_2_42
-- reg_a = a2_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001001000011",
--  (808) multiplication_with_reduction_special_prime_2_43
-- reg_a = o2_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001001010111",
--  (809) multiplication_with_reduction_special_prime_2_44
-- reg_a = a3_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
"001011100001100000000000100000000000000100000101100011",
--  (810) multiplication_with_reduction_special_prime_2_45
-- In case of size 5
-- reg_a = a0_X; reg_b = b4_X; reg_acc = reg_o; Enable sign b; operation : a*b + acc;
"000000100001100000000000100000000001000100010000000011",
--  (811) multiplication_with_reduction_special_prime_2_46
-- reg_a = a4_X; reg_b = b0_X; reg_acc = reg_o; o4_X = reg_o; Enable sign a; operation : a*b + acc;
"000000100001100000010000100000000000100010000010000011",
--  (812) multiplication_with_reduction_special_prime_2_47
-- reg_a = a1_X; reg_b = b4_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001100000000000100000100001000100010000100011",
--  (813) multiplication_with_reduction_special_prime_2_48
-- reg_a = o1_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100010000110111",
--  (814) multiplication_with_reduction_special_prime_2_49
-- reg_a = a2_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001101000011",
--  (815) multiplication_with_reduction_special_prime_2_50
-- reg_a = o2_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001101010111",
--  (816) multiplication_with_reduction_special_prime_2_51
-- reg_a = a3_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001001100011",
--  (817) multiplication_with_reduction_special_prime_2_52
-- reg_a = o3_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001001110111",
--  (818) multiplication_with_reduction_special_prime_2_53
-- reg_a = a4_X; reg_b = b1_X; reg_acc = reg_o; o0_X = reg_o; Enable sign a; operation : a*b + acc;
"000000100001100000010000100000000000100100000110000011",
--  (819) multiplication_with_reduction_special_prime_2_54
-- reg_a = a2_X; reg_b = b4_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001100000000000100000100001000100010001000011",
--  (820) multiplication_with_reduction_special_prime_2_55
-- reg_a = o2_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100010001010111",
--  (821) multiplication_with_reduction_special_prime_2_56
-- reg_a = a3_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001101100011",
--  (822) multiplication_with_reduction_special_prime_2_57
-- reg_a = o3_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001101110111",
--  (823) multiplication_with_reduction_special_prime_2_58
-- reg_a = a4_X; reg_b = b2_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001100000000000100000000000100100001010000011",
--  (824) multiplication_with_reduction_special_prime_2_59
-- reg_a = o4_X; reg_b = primeSP2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
"000000100001100000010000100000000000001000101010010111",
--  (825) multiplication_with_reduction_special_prime_2_60
-- reg_a = a3_X; reg_b = b4_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001100000000000100000100001000100010001100011",
--  (826) multiplication_with_reduction_special_prime_2_61
-- reg_a = o3_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100010001110111",
--  (827) multiplication_with_reduction_special_prime_2_62
-- reg_a = a4_X; reg_b = b3_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001100000000000100000000000100100001110000011",
--  (828) multiplication_with_reduction_special_prime_2_63
-- reg_a = o4_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
"000000100001100000010000100000000000001101001110010111",
--  (829) multiplication_with_reduction_special_prime_2_64
-- reg_a = a4_X; reg_b = b4_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001100000000000100000100001100100010010000011",
--  (830) multiplication_with_reduction_special_prime_2_65
-- reg_a = o4_X; reg_b = primeSP4; reg_acc = reg_o; o3_X = reg_o; o4_X = reg_o >> 256; operation : a*b + acc;
"000000100001100001110000100000000000010001110010010111",
--  (831) multiplication_with_reduction_special_prime_2_66
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (832) multiplication_with_reduction_special_prime_2_67
-- -- In case of sizes 6, 7, 8
-- reg_a = a0_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010000000011",
--  (833) multiplication_with_reduction_special_prime_2_68
-- reg_a = a4_X; reg_b = b0_X; reg_acc = reg_o; o4_X = reg_o; operation : a*b + acc;
"000000100001101000010000100000000000010010000010000011",
--  (834) multiplication_with_reduction_special_prime_2_69
-- reg_a = o0_X; reg_b = primeSP5; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001101000000000100000100000000100010100010111",
--  (835) multiplication_with_reduction_special_prime_2_70
-- reg_a = a1_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010000100011",
--  (836) multiplication_with_reduction_special_prime_2_71
-- reg_a = o1_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010000110111",
--  (837) multiplication_with_reduction_special_prime_2_72
-- reg_a = a2_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001101000011",
--  (838) multiplication_with_reduction_special_prime_2_73
-- reg_a = o2_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001101010111",
--  (839) multiplication_with_reduction_special_prime_2_74
-- reg_a = a3_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001001100011",
--  (840) multiplication_with_reduction_special_prime_2_75
-- reg_a = o3_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001001110111",
--  (841) multiplication_with_reduction_special_prime_2_76
-- reg_a = a4_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
"010000100001101000000000100000000000000100000110000011",
--  (842) multiplication_with_reduction_special_prime_2_77
-- In case of size 6
-- reg_a = a0_X; reg_b = b5_X; reg_acc = reg_o; Enable sign b; operation : a*b + acc;
"000000100001101000000000100000000001000100010100000011",
--  (843) multiplication_with_reduction_special_prime_2_78
-- reg_a = a5_X; reg_b = b0_X; reg_acc = reg_o; o5_X = reg_o; Enable sign a; operation : a*b + acc;
"000000100001101000010000100000000000100010100010100011",
--  (844) multiplication_with_reduction_special_prime_2_79
-- reg_a = a1_X; reg_b = b5_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001101000000000100000100001000100010100100011",
--  (845) multiplication_with_reduction_special_prime_2_80
-- reg_a = o1_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010100110111",
--  (846) multiplication_with_reduction_special_prime_2_81
-- reg_a = a2_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010001000011",
--  (847) multiplication_with_reduction_special_prime_2_82
-- reg_a = o2_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010001010111",
--  (848) multiplication_with_reduction_special_prime_2_83
-- reg_a = a3_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001101100011",
--  (849) multiplication_with_reduction_special_prime_2_84
-- reg_a = o3_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001101110111",
--  (850) multiplication_with_reduction_special_prime_2_85
-- reg_a = a4_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001010000011",
--  (851) multiplication_with_reduction_special_prime_2_86
-- reg_a = o4_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001010010111",
--  (852) multiplication_with_reduction_special_prime_2_87
-- reg_a = a5_X; reg_b = b1_X; reg_acc = reg_o; o0_X = reg_o; Enable sign a; operation : a*b + acc;
"000000100001101000010000100000000000100100000110100011",
--  (853) multiplication_with_reduction_special_prime_2_88
-- reg_a = a2_X; reg_b = b5_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001101000000000100000100001000100010101000011",
--  (854) multiplication_with_reduction_special_prime_2_89
-- reg_a = o2_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010101010111",
--  (855) multiplication_with_reduction_special_prime_2_90
-- reg_a = a3_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010001100011",
--  (856) multiplication_with_reduction_special_prime_2_91
-- reg_a = o3_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010001110111",
--  (857) multiplication_with_reduction_special_prime_2_92
-- reg_a = a4_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001110000011",
--  (858) multiplication_with_reduction_special_prime_2_93
-- reg_a = o4_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001110010111",
--  (859) multiplication_with_reduction_special_prime_2_94
-- reg_a = a5_X; reg_b = b2_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001101000000000100000000000100100001010100011",
--  (860) multiplication_with_reduction_special_prime_2_95
-- reg_a = o5_X; reg_b = primeSP2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
"000000100001101000010000100000000000001000101010110111",
--  (861) multiplication_with_reduction_special_prime_2_96
-- reg_a = a3_X; reg_b = b5_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001101000000000100000100001000100010101100011",
--  (862) multiplication_with_reduction_special_prime_2_97
-- reg_a = o3_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010101110111",
--  (863) multiplication_with_reduction_special_prime_2_98
-- reg_a = a4_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010010000011",
--  (864) multiplication_with_reduction_special_prime_2_99
-- reg_a = o4_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010010010111",
--  (865) multiplication_with_reduction_special_prime_2_100
-- reg_a = a5_X; reg_b = b3_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001101000000000100000000000100100001110100011",
--  (866) multiplication_with_reduction_special_prime_2_101
-- reg_a = o5_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
"000000100001101000010000100000000000001101001110110111",
--  (867) multiplication_with_reduction_special_prime_2_102
-- reg_a = a4_X; reg_b = b5_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001101000000000100000100001000100010110000011",
--  (868) multiplication_with_reduction_special_prime_2_103
-- reg_a = o4_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010110010111",
--  (869) multiplication_with_reduction_special_prime_2_104
-- reg_a = a5_X; reg_b = b4_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001101000000000100000000000100100010010100011",
--  (870) multiplication_with_reduction_special_prime_2_105
-- reg_a = o5_X; reg_b = primeSP4; reg_acc = reg_o; o3_X = reg_o; operation : a*b + acc;
"000000100001101000010000100000000000010001110010110111",
--  (871) multiplication_with_reduction_special_prime_2_106
-- reg_a = a5_X; reg_b = b5_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001101000000000100000100001100100010110100011",
--  (872) multiplication_with_reduction_special_prime_2_107
-- reg_a = o5_X; reg_b = primeSP5; reg_acc = reg_o; o4_X = reg_o; o5_X = reg_o >> 256; operation : a*b + acc;
"000000100001101001110000100000000000010110010110110111",
--  (873) multiplication_with_reduction_special_prime_2_108
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (874) multiplication_with_reduction_special_prime_2_109
-- -- In case of sizes 7, 8
-- reg_a = a0_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010100000011",
--  (875) multiplication_with_reduction_special_prime_2_110
-- reg_a = a5_X; reg_b = b0_X; reg_acc = reg_o; o5_X = reg_o; operation : a*b + acc;
"000000100001110000010000100000000000011010100010100011",
--  (876) multiplication_with_reduction_special_prime_2_111
-- reg_a = o0_X; reg_b = primeSP6; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001110000000000100000100000000100011000010111",
--  (877) multiplication_with_reduction_special_prime_2_112
-- reg_a = a1_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010100100011",
--  (878) multiplication_with_reduction_special_prime_2_113
-- reg_a = o1_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010100110111",
--  (879) multiplication_with_reduction_special_prime_2_114
-- reg_a = a2_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010001000011",
--  (880) multiplication_with_reduction_special_prime_2_115
-- reg_a = o2_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010001010111",
--  (881) multiplication_with_reduction_special_prime_2_116
-- reg_a = a3_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001101100011",
--  (882) multiplication_with_reduction_special_prime_2_117
-- reg_a = o3_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001101110111",
--  (883) multiplication_with_reduction_special_prime_2_118
-- reg_a = a4_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001010000011",
--  (884) multiplication_with_reduction_special_prime_2_119
-- reg_a = o4_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001010010111",
--  (885) multiplication_with_reduction_special_prime_2_120
-- reg_a = a5_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
"010110100001110000000000100000000000000100000110100011",
--  (886) multiplication_with_reduction_special_prime_2_121
-- -- In case of size 7
-- reg_a = a0_X; reg_b = b6_X; reg_acc = reg_o; Enable sign b; operation : a*b + acc;
"000000100001110000000000100000000001000100011000000011",
--  (887) multiplication_with_reduction_special_prime_2_122
-- reg_a = a6_X; reg_b = b0_X; reg_acc = reg_o; o6_X = reg_o; Enable sign a; operation : a*b + acc;
"000000100001110000010000100000000000100011000011000011",
--  (888) multiplication_with_reduction_special_prime_2_123
-- reg_a = a1_X; reg_b = b6_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001110000000000100000100001000100011000100011",
--  (889) multiplication_with_reduction_special_prime_2_124
-- reg_a = o1_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100011000110111",
--  (890) multiplication_with_reduction_special_prime_2_125
-- reg_a = a2_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010101000011",
--  (891) multiplication_with_reduction_special_prime_2_126
-- reg_a = o2_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010101010111",
--  (892) multiplication_with_reduction_special_prime_2_127
-- reg_a = a3_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010001100011",
--  (893) multiplication_with_reduction_special_prime_2_128
-- reg_a = o3_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010001110111",
--  (894) multiplication_with_reduction_special_prime_2_129
-- reg_a = a4_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001110000011",
--  (895) multiplication_with_reduction_special_prime_2_130
-- reg_a = o4_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001110010111",
--  (896) multiplication_with_reduction_special_prime_2_131
-- reg_a = a5_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001010100011",
--  (897) multiplication_with_reduction_special_prime_2_132
-- reg_a = o5_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001010110111",
--  (898) multiplication_with_reduction_special_prime_2_133
-- reg_a = a6_X; reg_b = b1_X; reg_acc = reg_o; Enable sign a; o0_X = reg_o; operation : a*b + acc;
"000000100001110000010000100000000000100100000111000011",
--  (899) multiplication_with_reduction_special_prime_2_134
-- reg_a = a2_X; reg_b = b6_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001110000000000100000100001000100011001000011",
--  (900) multiplication_with_reduction_special_prime_2_135
-- reg_a = o2_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100011001010111",
--  (901) multiplication_with_reduction_special_prime_2_136
-- reg_a = a3_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010101100011",
--  (902) multiplication_with_reduction_special_prime_2_137
-- reg_a = o3_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010101110111",
--  (903) multiplication_with_reduction_special_prime_2_138
-- reg_a = a4_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010010000011",
--  (904) multiplication_with_reduction_special_prime_2_139
-- reg_a = o4_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010010010111",
--  (905) multiplication_with_reduction_special_prime_2_140
-- reg_a = a5_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001110100011",
--  (906) multiplication_with_reduction_special_prime_2_141
-- reg_a = o5_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001110110111",
--  (907) multiplication_with_reduction_special_prime_2_142
-- reg_a = a6_X; reg_b = b2_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001110000000000100000000000100100001011000011",
--  (908) multiplication_with_reduction_special_prime_2_143
-- reg_a = o6_X; reg_b = primeSP2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
"000000100001110000010000100000000000001000101011010111",
--  (909) multiplication_with_reduction_special_prime_2_144
-- reg_a = a3_X; reg_b = b6_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001110000000000100000100001000100011001100011",
--  (910) multiplication_with_reduction_special_prime_2_145
-- reg_a = o3_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100011001110111",
--  (911) multiplication_with_reduction_special_prime_2_146
-- reg_a = a4_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010110000011",
--  (912) multiplication_with_reduction_special_prime_2_147
-- reg_a = o4_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010110010111",
--  (913) multiplication_with_reduction_special_prime_2_148
-- reg_a = a5_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010010100011",
--  (914) multiplication_with_reduction_special_prime_2_149
-- reg_a = o5_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010010110111",
--  (915) multiplication_with_reduction_special_prime_2_150
-- reg_a = a6_X; reg_b = b3_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001110000000000100000000000100100001111000011",
--  (916) multiplication_with_reduction_special_prime_2_151
-- reg_a = o6_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
"000000100001110000010000100000000000001101001111010111",
--  (917) multiplication_with_reduction_special_prime_2_152
-- reg_a = a4_X; reg_b = b6_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001110000000000100000100001000100011010000011",
--  (918) multiplication_with_reduction_special_prime_2_153
-- reg_a = o4_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100011010010111",
--  (919) multiplication_with_reduction_special_prime_2_154
-- reg_a = a5_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010110100011",
--  (920) multiplication_with_reduction_special_prime_2_155
-- reg_a = o5_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010110110111",
--  (921) multiplication_with_reduction_special_prime_2_156
-- reg_a = a6_X; reg_b = b4_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001110000000000100000000000100100010011000011",
--  (922) multiplication_with_reduction_special_prime_2_157
-- reg_a = o6_X; reg_b = primeSP4; reg_acc = reg_o; o3_X = reg_o; operation : a*b + acc;
"000000100001110000010000100000000000010001110011010111",
--  (923) multiplication_with_reduction_special_prime_2_158
-- reg_a = a5_X; reg_b = b6_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001110000000000100000100001000100011010100011",
--  (924) multiplication_with_reduction_special_prime_2_159
-- reg_a = o5_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100011010110111",
--  (925) multiplication_with_reduction_special_prime_2_160
-- reg_a = a6_X; reg_b = b5_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001110000000000100000000000100100010111000011",
--  (926) multiplication_with_reduction_special_prime_2_161
-- reg_a = o6_X; reg_b = primeSP5; reg_acc = reg_o; o4_X = reg_o; operation : a*b + acc;
"000000100001110000010000100000000000010110010111010111",
--  (927) multiplication_with_reduction_special_prime_2_162
-- reg_a = a6_X; reg_b = b6_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001110000000000100000100001100100011011000011",
--  (928) multiplication_with_reduction_special_prime_2_163
-- reg_a = o6_X; reg_b = primeSP6; reg_acc = reg_o; o5_X = reg_o; o6_X = reg_o >> 256; operation : a*b + acc;
"000000100001110001110000100000000000011010111011010111",
--  (929) multiplication_with_reduction_special_prime_2_164
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (930) multiplication_with_reduction_special_prime_2_165
-- -- In case of size 8
-- reg_a = a0_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011000000011",
--  (931) multiplication_with_reduction_special_prime_2_166
-- reg_a = a6_X; reg_b = b0_X; reg_acc = reg_o; o6_X = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000011011000011000011",
--  (932) multiplication_with_reduction_special_prime_2_167
-- reg_a = o0_X; reg_b = primeSP7; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001111000000000100000100000000100011100010111",
--  (933) multiplication_with_reduction_special_prime_2_168
-- reg_a = a1_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011000100011",
--  (934) multiplication_with_reduction_special_prime_2_169
-- reg_a = o1_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011000110111",
--  (935) multiplication_with_reduction_special_prime_2_170
-- reg_a = a2_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010101000011",
--  (936) multiplication_with_reduction_special_prime_2_171
-- reg_a = o2_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010101010111",
--  (937) multiplication_with_reduction_special_prime_2_172
-- reg_a = a3_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010001100011",
--  (938) multiplication_with_reduction_special_prime_2_173
-- reg_a = o3_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010001110111",
--  (939) multiplication_with_reduction_special_prime_2_174
-- reg_a = a4_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001110000011",
--  (940) multiplication_with_reduction_special_prime_2_175
-- reg_a = o4_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001110010111",
--  (941) multiplication_with_reduction_special_prime_2_176
-- reg_a = a5_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001010100011",
--  (942) multiplication_with_reduction_special_prime_2_177
-- reg_a = o5_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001010110111",
--  (943) multiplication_with_reduction_special_prime_2_178
-- reg_a = a6_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100000111000011",
--  (944) multiplication_with_reduction_special_prime_2_179
-- reg_a = a0_X; reg_b = b7_X; reg_acc = reg_o; Enable sign b; operation : a*b + acc;
"000000100001111000000000100000000001000100011100000011",
--  (945) multiplication_with_reduction_special_prime_2_180
-- reg_a = a7_X; reg_b = b0_X; reg_acc = reg_o; o7_X = reg_o; Enable sign a; operation : a*b + acc;
"000000100001111000010000100000000000100011100011100011",
--  (946) multiplication_with_reduction_special_prime_2_181
-- reg_a = a1_X; reg_b = b7_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001111000000000100000100001000100011100100011",
--  (947) multiplication_with_reduction_special_prime_2_182
-- reg_a = o1_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011100110111",
--  (948) multiplication_with_reduction_special_prime_2_183
-- reg_a = a2_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011001000011",
--  (949) multiplication_with_reduction_special_prime_2_184
-- reg_a = o2_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011001010111",
--  (950) multiplication_with_reduction_special_prime_2_185
-- reg_a = a3_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010101100011",
--  (951) multiplication_with_reduction_special_prime_2_186
-- reg_a = o3_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010101110111",
--  (952) multiplication_with_reduction_special_prime_2_187
-- reg_a = a4_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010010000011",
--  (953) multiplication_with_reduction_special_prime_2_188
-- reg_a = o4_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010010010111",
--  (954) multiplication_with_reduction_special_prime_2_189
-- reg_a = a5_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001110100011",
--  (955) multiplication_with_reduction_special_prime_2_190
-- reg_a = o5_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001110110111",
--  (956) multiplication_with_reduction_special_prime_2_191
-- reg_a = a6_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001011000011",
--  (957) multiplication_with_reduction_special_prime_2_192
-- reg_a = o6_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001011010111",
--  (958) multiplication_with_reduction_special_prime_2_193
-- reg_a = a7_X; reg_b = b1_X; reg_acc = reg_o; Enable sign a; o0_X = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000100100000111100011",
--  (959) multiplication_with_reduction_special_prime_2_194
-- reg_a = a2_X; reg_b = b7_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001111000000000100000100001000100011101000011",
--  (960) multiplication_with_reduction_special_prime_2_195
-- reg_a = o2_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011101010111",
--  (961) multiplication_with_reduction_special_prime_2_196
-- reg_a = a3_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011001100011",
--  (962) multiplication_with_reduction_special_prime_2_197
-- reg_a = o3_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011001110111",
--  (963) multiplication_with_reduction_special_prime_2_198
-- reg_a = a4_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010110000011",
--  (964) multiplication_with_reduction_special_prime_2_199
-- reg_a = o4_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010110010111",
--  (965) multiplication_with_reduction_special_prime_2_200
-- reg_a = a5_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010010100011",
--  (966) multiplication_with_reduction_special_prime_2_201
-- reg_a = o5_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010010110111",
--  (967) multiplication_with_reduction_special_prime_2_202
-- reg_a = a6_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001111000011",
--  (968) multiplication_with_reduction_special_prime_2_203
-- reg_a = o6_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001111010111",
--  (969) multiplication_with_reduction_special_prime_2_204
-- reg_a = a7_X; reg_b = b2_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001111000000000100000000000100100001011100011",
--  (970) multiplication_with_reduction_special_prime_2_205
-- reg_a = o7_X; reg_b = primeSP2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000001000101011110111",
--  (971) multiplication_with_reduction_special_prime_2_206
-- reg_a = a3_X; reg_b = b7_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001111000000000100000100001000100011101100011",
--  (972) multiplication_with_reduction_special_prime_2_207
-- reg_a = o3_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011101110111",
--  (973) multiplication_with_reduction_special_prime_2_208
-- reg_a = a4_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011010000011",
--  (974) multiplication_with_reduction_special_prime_2_209
-- reg_a = o4_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011010010111",
--  (975) multiplication_with_reduction_special_prime_2_210
-- reg_a = a5_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010110100011",
--  (976) multiplication_with_reduction_special_prime_2_211
-- reg_a = o5_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010110110111",
--  (977) multiplication_with_reduction_special_prime_2_212
-- reg_a = a6_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010011000011",
--  (978) multiplication_with_reduction_special_prime_2_213
-- reg_a = o6_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010011010111",
--  (979) multiplication_with_reduction_special_prime_2_214
-- reg_a = a7_X; reg_b = b3_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001111000000000100000000000100100001111100011",
--  (980) multiplication_with_reduction_special_prime_2_215
-- reg_a = o7_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000001101001111110111",
--  (981) multiplication_with_reduction_special_prime_2_216
-- reg_a = a4_X; reg_b = b7_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001111000000000100000100001000100011110000011",
--  (982) multiplication_with_reduction_special_prime_2_217
-- reg_a = o4_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011110010111",
--  (983) multiplication_with_reduction_special_prime_2_218
-- reg_a = a5_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011010100011",
--  (984) multiplication_with_reduction_special_prime_2_219
-- reg_a = o5_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011010110111",
--  (985) multiplication_with_reduction_special_prime_2_220
-- reg_a = a6_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010111000011",
--  (986) multiplication_with_reduction_special_prime_2_221
-- reg_a = o6_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010111010111",
--  (987) multiplication_with_reduction_special_prime_2_222
-- reg_a = a7_X; reg_b = b4_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001111000000000100000000000100100010011100011",
--  (988) multiplication_with_reduction_special_prime_2_223
-- reg_a = o7_X; reg_b = primeSP4; reg_acc = reg_o; o3_X = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000010001110011110111",
--  (989) multiplication_with_reduction_special_prime_2_224
-- reg_a = a5_X; reg_b = b7_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001111000000000100000100001000100011110100011",
--  (990) multiplication_with_reduction_special_prime_2_225
-- reg_a = o5_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011110110111",
--  (991) multiplication_with_reduction_special_prime_2_226
-- reg_a = a6_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011011000011",
--  (992) multiplication_with_reduction_special_prime_2_227
-- reg_a = o6_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011011010111",
--  (993) multiplication_with_reduction_special_prime_2_228
-- reg_a = a7_X; reg_b = b5_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001111000000000100000000000100100010111100011",
--  (994) multiplication_with_reduction_special_prime_2_229
-- reg_a = o7_X; reg_b = primeSP5; reg_acc = reg_o; o4_X = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000010110010111110111",
--  (995) multiplication_with_reduction_special_prime_2_230
-- reg_a = a6_X; reg_b = b7_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001111000000000100000100001000100011111000011",
--  (996) multiplication_with_reduction_special_prime_2_231
-- reg_a = o6_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011111010111",
--  (997) multiplication_with_reduction_special_prime_2_232
-- reg_a = a7_X; reg_b = b6_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001111000000000100000000000100100011011100011",
--  (998) multiplication_with_reduction_special_prime_2_233
-- reg_a = o7_X; reg_b = primeSP6; reg_acc = reg_o; o5_X = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000011010111011110111",
--  (999) multiplication_with_reduction_special_prime_2_234
-- reg_a = a7_X; reg_b = b7_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001111000000000100000100001100100011111100011",
--  (1000) multiplication_with_reduction_special_prime_2_235
-- reg_a = o7_X; reg_b = primeSP7; reg_acc = reg_o; o6_X = reg_o; o7_X = reg_o >> 256; operation : a*b + acc;
"000000100001111001110000100000000000011111011111110111",
--  (1001) multiplication_with_reduction_special_prime_2_236
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (1002) multiplication_with_reduction_special_prime_3_0
-- -- In case of sizes 3, 4, 5, 6, 7, 8
-- reg_a = a0_X; reg_b = b0_X; reg_acc = 0; o0_X = reg_o; operation : a*b + acc;
"000000100001010000010000100000010000000100000000000011",
--  (1003) multiplication_with_reduction_special_prime_3_1
-- reg_a = a0_X; reg_b = b1_X; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001010000000000100000100000000100000100000011",
--  (1004) multiplication_with_reduction_special_prime_3_2
-- reg_a = a1_X; reg_b = b0_X; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
"000000100001010000010000100000000000001000100000100011",
--  (1005) multiplication_with_reduction_special_prime_3_3
-- reg_a = a1_X; reg_b = b1_X; reg_acc = reg_o >> 256; operation : a*b + acc;
"000011100001010000000000100000100000000100000100100011",
--  (1006) multiplication_with_reduction_special_prime_3_4
-- -- In case of size 3
-- reg_a = a0_X; reg_b = b2_X; reg_acc = reg_o; Enable sign b; operation : a*b + acc;
"000000100001010000000000100000000001000100001000000011",
--  (1007) multiplication_with_reduction_special_prime_3_5
-- reg_a = a2_X; reg_b = b0_X; reg_acc = reg_o; o2_X = reg_o; Enable sign a; operation : a*b + acc;
"000000100001010000010000100000000000101101000001000011",
--  (1008) multiplication_with_reduction_special_prime_3_6
-- reg_a = a1_X; reg_b = b2_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001010000000000100000100001000100001000100011",
--  (1009) multiplication_with_reduction_special_prime_3_7
-- reg_a = a2_X; reg_b = b1_X; reg_acc = reg_o; Enable sign a; o0_X = reg_o; operation : a*b + acc;
"000000100001010000010000100000000000100100000101000011",
--  (1010) multiplication_with_reduction_special_prime_3_8
-- reg_a = a2_X; reg_b = b2_X; reg_acc = reg_o >> 256; Enable sign a,b; o1_X = reg_o; o2_X = reg_o >> 256; operation : a*b + acc;
"000000100001010001110000100000100001100100001001000011",
--  (1011) multiplication_with_reduction_special_prime_3_9
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (1012) multiplication_with_reduction_special_prime_3_10
-- -- In case of sizes 4, 5, 6, 7, 8
-- reg_a = a0_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001011000000000100000000000000100001000000011",
--  (1013) multiplication_with_reduction_special_prime_3_11
-- reg_a = a2_X; reg_b = b0_X; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
"000000100001011000010000100000000000001101000001000011",
--  (1014) multiplication_with_reduction_special_prime_3_12
-- reg_a = o0_X; reg_b = primeSP3; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001011000000000100000100000000100001100010111",
--  (1015) multiplication_with_reduction_special_prime_3_13
-- reg_a = a1_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001011000000000100000000000000100001000100011",
--  (1016) multiplication_with_reduction_special_prime_3_14
-- reg_a = a2_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
"000110100001011000000000100000000000000100000101000011",
--  (1017) multiplication_with_reduction_special_prime_3_15
-- -- In case of size 4
-- reg_a = a0_X; reg_b = b3_X; reg_acc = reg_o; Enable sign b; operation : a*b + acc;
"000000100001011000000000100000000001000100001100000011",
--  (1018) multiplication_with_reduction_special_prime_3_16
-- reg_a = a3_X; reg_b = b0_X; reg_acc = reg_o; o3_X = reg_o; Enable sign a; operation : a*b + acc;
"000000100001011000010000100000000000100001100001100011",
--  (1019) multiplication_with_reduction_special_prime_3_17
-- reg_a = a1_X; reg_b = b3_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001011000000000100000100001000100001100100011",
--  (1020) multiplication_with_reduction_special_prime_3_18
-- reg_a = o1_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001011000000000100000000000000100001100110111",
--  (1021) multiplication_with_reduction_special_prime_3_19
-- reg_a = a2_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001011000000000100000000000000100001001000011",
--  (1022) multiplication_with_reduction_special_prime_3_20
-- reg_a = a3_X; reg_b = b1_X; reg_acc = reg_o; Enable sign a; o0_X = reg_o; operation : a*b + acc;
"000000100001011000010000100000000000100100000101100011",
--  (1023) multiplication_with_reduction_special_prime_3_21
-- reg_a = a2_X; reg_b = b3_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001011000000000100000100001000100001101000011",
--  (1024) multiplication_with_reduction_special_prime_3_22
-- reg_a = o2_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001011000000000100000000000000100001101010111",
--  (1025) multiplication_with_reduction_special_prime_3_23
-- reg_a = a3_X; reg_b = b2_X; reg_acc = reg_o; Enable sign a; o1_X = reg_o; operation : a*b + acc;
"000000100001011000010000100000000000101000101001100011",
--  (1026) multiplication_with_reduction_special_prime_3_24
-- reg_a = a3_X; reg_b = b3_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001011000000000100000100001100100001101100011",
--  (1027) multiplication_with_reduction_special_prime_3_25
-- reg_a = o3_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; o3_X = reg_o >> 256; operation : a*b + acc;
"000000100001011001110000100000000000001101001101110111",
--  (1028) multiplication_with_reduction_special_prime_3_26
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (1029) multiplication_with_reduction_special_prime_3_27
-- -- In case of sizes 5, 6, 7, 8
-- reg_a = a0_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001100000011",
--  (1030) multiplication_with_reduction_special_prime_3_28
-- reg_a = a3_X; reg_b = b0_X; reg_acc = reg_o; o3_X = reg_o; operation : a*b + acc;
"000000100001100000010000100000000000010001100001100011",
--  (1031) multiplication_with_reduction_special_prime_3_29
-- reg_a = o0_X; reg_b = primeSP4; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001100000000000100000100000000100010000010111",
--  (1032) multiplication_with_reduction_special_prime_3_30
-- reg_a = a1_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001100100011",
--  (1033) multiplication_with_reduction_special_prime_3_31
-- reg_a = o1_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001100110111",
--  (1034) multiplication_with_reduction_special_prime_3_32
-- reg_a = a2_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001001000011",
--  (1035) multiplication_with_reduction_special_prime_3_33
-- reg_a = a3_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
"001010100001100000000000100000000000000100000101100011",
--  (1036) multiplication_with_reduction_special_prime_3_34
-- In case of size 5
-- reg_a = a0_X; reg_b = b4_X; reg_acc = reg_o; Enable sign b; operation : a*b + acc;
"000000100001100000000000100000000001000100010000000011",
--  (1037) multiplication_with_reduction_special_prime_3_35
-- reg_a = a4_X; reg_b = b0_X; reg_acc = reg_o; o4_X = reg_o; Enable sign a; operation : a*b + acc;
"000000100001100000010000100000000000100010000010000011",
--  (1038) multiplication_with_reduction_special_prime_3_36
-- reg_a = a1_X; reg_b = b4_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001100000000000100000100001000100010000100011",
--  (1039) multiplication_with_reduction_special_prime_3_37
-- reg_a = o1_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100010000110111",
--  (1040) multiplication_with_reduction_special_prime_3_38
-- reg_a = a2_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001101000011",
--  (1041) multiplication_with_reduction_special_prime_3_39
-- reg_a = o2_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001101010111",
--  (1042) multiplication_with_reduction_special_prime_3_40
-- reg_a = a3_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001001100011",
--  (1043) multiplication_with_reduction_special_prime_3_41
-- reg_a = a4_X; reg_b = b1_X; reg_acc = reg_o; o0_X = reg_o; Enable sign a; operation : a*b + acc;
"000000100001100000010000100000000000100100000110000011",
--  (1044) multiplication_with_reduction_special_prime_3_42
-- reg_a = a2_X; reg_b = b4_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001100000000000100000100001000100010001000011",
--  (1045) multiplication_with_reduction_special_prime_3_43
-- reg_a = o2_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100010001010111",
--  (1046) multiplication_with_reduction_special_prime_3_44
-- reg_a = a3_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001101100011",
--  (1047) multiplication_with_reduction_special_prime_3_45
-- reg_a = o3_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001101110111",
--  (1048) multiplication_with_reduction_special_prime_3_46
-- reg_a = a4_X; reg_b = b2_X; reg_acc = reg_o; Enable sign a; o1_X = reg_o; operation : a*b + acc;
"000000100001100000010000100000000000101000101010000011",
--  (1049) multiplication_with_reduction_special_prime_3_47
-- reg_a = a3_X; reg_b = b4_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001100000000000100000100001000100010001100011",
--  (1050) multiplication_with_reduction_special_prime_3_48
-- reg_a = o3_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100010001110111",
--  (1051) multiplication_with_reduction_special_prime_3_49
-- reg_a = a4_X; reg_b = b3_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001100000000000100000000000100100001110000011",
--  (1052) multiplication_with_reduction_special_prime_3_50
-- reg_a = o4_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
"000000100001100000010000100000000000001101001110010111",
--  (1053) multiplication_with_reduction_special_prime_3_51
-- reg_a = a4_X; reg_b = b4_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001100000000000100000100001100100010010000011",
--  (1054) multiplication_with_reduction_special_prime_3_52
-- reg_a = o4_X; reg_b = primeSP4; reg_acc = reg_o; o3_X = reg_o; o4_X = reg_o >> 256; operation : a*b + acc;
"000000100001100001110000100000000000010001110010010111",
--  (1055) multiplication_with_reduction_special_prime_3_53
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (1056) multiplication_with_reduction_special_prime_3_54
-- -- In case of sizes 6, 7, 8
-- reg_a = a0_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010000000011",
--  (1057) multiplication_with_reduction_special_prime_3_55
-- reg_a = a4_X; reg_b = b0_X; reg_acc = reg_o; o4_X = reg_o; operation : a*b + acc;
"000000100001101000010000100000000000010110000010000011",
--  (1058) multiplication_with_reduction_special_prime_3_56
-- reg_a = o0_X; reg_b = primeSP5; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001101000000000100000100000000100010100010111",
--  (1059) multiplication_with_reduction_special_prime_3_57
-- reg_a = a1_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010000100011",
--  (1060) multiplication_with_reduction_special_prime_3_58
-- reg_a = o1_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010000110111",
--  (1061) multiplication_with_reduction_special_prime_3_59
-- reg_a = a2_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001101000011",
--  (1062) multiplication_with_reduction_special_prime_3_60
-- reg_a = o2_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001101010111",
--  (1063) multiplication_with_reduction_special_prime_3_61
-- reg_a = a3_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001001100011",
--  (1064) multiplication_with_reduction_special_prime_3_62
-- reg_a = a4_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
"001111100001101000000000100000000000000100000110000011",
--  (1065) multiplication_with_reduction_special_prime_3_63
-- In case of size 6
-- reg_a = a0_X; reg_b = b5_X; reg_acc = reg_o; Enable sign b; operation : a*b + acc;
"000000100001101000000000100000000001000100010100000011",
--  (1066) multiplication_with_reduction_special_prime_3_64
-- reg_a = a5_X; reg_b = b0_X; reg_acc = reg_o; o5_X = reg_o; Enable sign a; operation : a*b + acc;
"000000100001101000010000100000000000100010100010100011",
--  (1067) multiplication_with_reduction_special_prime_3_65
-- reg_a = a1_X; reg_b = b5_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001101000000000100000100001000100010100100011",
--  (1068) multiplication_with_reduction_special_prime_3_66
-- reg_a = o1_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010100110111",
--  (1069) multiplication_with_reduction_special_prime_3_67
-- reg_a = a2_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010001000011",
--  (1070) multiplication_with_reduction_special_prime_3_68
-- reg_a = o2_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010001010111",
--  (1071) multiplication_with_reduction_special_prime_3_69
-- reg_a = a3_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001101100011",
--  (1072) multiplication_with_reduction_special_prime_3_70
-- reg_a = o3_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001101110111",
--  (1073) multiplication_with_reduction_special_prime_3_71
-- reg_a = a4_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001010000011",
--  (1074) multiplication_with_reduction_special_prime_3_72
-- reg_a = a5_X; reg_b = b1_X; reg_acc = reg_o; o0_X = reg_o; Enable sign a; operation : a*b + acc;
"000000100001101000010000100000000000100100000110100011",
--  (1075) multiplication_with_reduction_special_prime_3_73
-- reg_a = a2_X; reg_b = b5_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001101000000000100000100001000100010101000011",
--  (1076) multiplication_with_reduction_special_prime_3_74
-- reg_a = o2_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010101010111",
--  (1077) multiplication_with_reduction_special_prime_3_75
-- reg_a = a3_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010001100011",
--  (1078) multiplication_with_reduction_special_prime_3_76
-- reg_a = o3_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010001110111",
--  (1079) multiplication_with_reduction_special_prime_3_77
-- reg_a = a4_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001110000011",
--  (1080) multiplication_with_reduction_special_prime_3_78
-- reg_a = o4_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001110010111",
--  (1081) multiplication_with_reduction_special_prime_3_79
-- reg_a = a5_X; reg_b = b2_X; reg_acc = reg_o; Enable sign a; o1_X = reg_o; operation : a*b + acc;
"000000100001101000010000100000000000101000101010100011",
--  (1082) multiplication_with_reduction_special_prime_3_80
-- reg_a = a3_X; reg_b = b5_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001101000000000100000100001000100010101100011",
--  (1083) multiplication_with_reduction_special_prime_3_81
-- reg_a = o3_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010101110111",
--  (1084) multiplication_with_reduction_special_prime_3_82
-- reg_a = a4_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010010000011",
--  (1085) multiplication_with_reduction_special_prime_3_83
-- reg_a = o4_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010010010111",
--  (1086) multiplication_with_reduction_special_prime_3_84
-- reg_a = a5_X; reg_b = b3_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001101000000000100000000000100100001110100011",
--  (1087) multiplication_with_reduction_special_prime_3_85
-- reg_a = o5_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
"000000100001101000010000100000000000001101001110110111",
--  (1088) multiplication_with_reduction_special_prime_3_86
-- reg_a = a4_X; reg_b = b5_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001101000000000100000100001000100010110000011",
--  (1089) multiplication_with_reduction_special_prime_3_87
-- reg_a = o4_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010110010111",
--  (1090) multiplication_with_reduction_special_prime_3_88
-- reg_a = a5_X; reg_b = b4_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001101000000000100000000000100100010010100011",
--  (1091) multiplication_with_reduction_special_prime_3_89
-- reg_a = o5_X; reg_b = primeSP4; reg_acc = reg_o; o3_X = reg_o; operation : a*b + acc;
"000000100001101000010000100000000000010001110010110111",
--  (1092) multiplication_with_reduction_special_prime_3_90
-- reg_a = a5_X; reg_b = b5_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001101000000000100000100001100100010110100011",
--  (1093) multiplication_with_reduction_special_prime_3_91
-- reg_a = o5_X; reg_b = primeSP5; reg_acc = reg_o; o4_X = reg_o; o5_X = reg_o >> 256; operation : a*b + acc;
"000000100001101001110000100000000000010110010110110111",
--  (1094) multiplication_with_reduction_special_prime_3_92
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (1095) multiplication_with_reduction_special_prime_3_93
-- -- In case of sizes 7, 8
-- reg_a = a0_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010100000011",
--  (1096) multiplication_with_reduction_special_prime_3_94
-- reg_a = a5_X; reg_b = b0_X; reg_acc = reg_o; o5_X = reg_o; operation : a*b + acc;
"000000100001110000010000100000000000011010100010100011",
--  (1097) multiplication_with_reduction_special_prime_3_95
-- reg_a = o0_X; reg_b = primeSP6; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001110000000000100000100000000100011000010111",
--  (1098) multiplication_with_reduction_special_prime_3_96
-- reg_a = a1_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010100100011",
--  (1099) multiplication_with_reduction_special_prime_3_97
-- reg_a = o1_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010100110111",
--  (1100) multiplication_with_reduction_special_prime_3_98
-- reg_a = a2_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010001000011",
--  (1101) multiplication_with_reduction_special_prime_3_99
-- reg_a = o2_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010001010111",
--  (1102) multiplication_with_reduction_special_prime_3_100
-- reg_a = a3_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001101100011",
--  (1103) multiplication_with_reduction_special_prime_3_101
-- reg_a = o3_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001101110111",
--  (1104) multiplication_with_reduction_special_prime_3_102
-- reg_a = a4_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001010000011",
--  (1105) multiplication_with_reduction_special_prime_3_103
-- reg_a = a5_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
"010101100001110000000000100000000000000100000110100011",
--  (1106) multiplication_with_reduction_special_prime_3_104
-- -- In case of size 7
-- reg_a = a0_X; reg_b = b6_X; reg_acc = reg_o; Enable sign b; operation : a*b + acc;
"000000100001110000000000100000000001000100011000000011",
--  (1107) multiplication_with_reduction_special_prime_3_105
-- reg_a = a6_X; reg_b = b0_X; reg_acc = reg_o; o6_X = reg_o; Enable sign a; operation : a*b + acc;
"000000100001110000010000100000000000111111000011000011",
--  (1108) multiplication_with_reduction_special_prime_3_106
-- reg_a = a1_X; reg_b = b6_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001110000000000100000100001000100011000100011",
--  (1109) multiplication_with_reduction_special_prime_3_107
-- reg_a = o1_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100011000110111",
--  (1110) multiplication_with_reduction_special_prime_3_108
-- reg_a = a2_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010101000011",
--  (1111) multiplication_with_reduction_special_prime_3_109
-- reg_a = o2_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010101010111",
--  (1112) multiplication_with_reduction_special_prime_3_110
-- reg_a = a3_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010001100011",
--  (1113) multiplication_with_reduction_special_prime_3_111
-- reg_a = o3_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010001110111",
--  (1114) multiplication_with_reduction_special_prime_3_112
-- reg_a = a4_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001110000011",
--  (1115) multiplication_with_reduction_special_prime_3_113
-- reg_a = o4_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001110010111",
--  (1116) multiplication_with_reduction_special_prime_3_114
-- reg_a = a5_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001010100011",
--  (1117) multiplication_with_reduction_special_prime_3_115
-- reg_a = a6_X; reg_b = b1_X; reg_acc = reg_o; o0_X = reg_o; Enable sign a; operation : a*b + acc;
"000000100001110000010000100000000000100100000111000011",
--  (1118) multiplication_with_reduction_special_prime_3_116
-- reg_a = a2_X; reg_b = b6_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001110000000000100000100001000100011001000011",
--  (1119) multiplication_with_reduction_special_prime_3_117
-- reg_a = o2_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100011001010111",
--  (1120) multiplication_with_reduction_special_prime_3_118
-- reg_a = a3_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010101100011",
--  (1121) multiplication_with_reduction_special_prime_3_119
-- reg_a = o3_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010101110111",
--  (1122) multiplication_with_reduction_special_prime_3_120
-- reg_a = a4_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010010000011",
--  (1123) multiplication_with_reduction_special_prime_3_121
-- reg_a = o4_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010010010111",
--  (1124) multiplication_with_reduction_special_prime_3_122
-- reg_a = a5_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001110100011",
--  (1125) multiplication_with_reduction_special_prime_3_123
-- reg_a = o5_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001110110111",
--  (1126) multiplication_with_reduction_special_prime_3_124
-- reg_a = a6_X; reg_b = b2_X; reg_acc = reg_o; o1_X = reg_o; Enable sign a; operation : a*b + acc;
"000000100001110000010000100000000000101000101011000011",
--  (1127) multiplication_with_reduction_special_prime_3_125
-- reg_a = a3_X; reg_b = b6_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001110000000000100000100001000100011001100011",
--  (1128) multiplication_with_reduction_special_prime_3_126
-- reg_a = o3_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100011001110111",
--  (1129) multiplication_with_reduction_special_prime_3_127
-- reg_a = a4_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010110000011",
--  (1130) multiplication_with_reduction_special_prime_3_128
-- reg_a = o4_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010110010111",
--  (1131) multiplication_with_reduction_special_prime_3_129
-- reg_a = a5_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010010100011",
--  (1132) multiplication_with_reduction_special_prime_3_130
-- reg_a = o5_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010010110111",
--  (1133) multiplication_with_reduction_special_prime_3_131
-- reg_a = a6_X; reg_b = b3_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001110000000000100000000000100100001111000011",
--  (1134) multiplication_with_reduction_special_prime_3_132
-- reg_a = o6_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
"000000100001110000010000100000000000001101001111010111",
--  (1135) multiplication_with_reduction_special_prime_3_133
-- reg_a = a4_X; reg_b = b6_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001110000000000100000100001000100011010000011",
--  (1136) multiplication_with_reduction_special_prime_3_134
-- reg_a = o4_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100011010010111",
--  (1137) multiplication_with_reduction_special_prime_3_135
-- reg_a = a5_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010110100011",
--  (1138) multiplication_with_reduction_special_prime_3_136
-- reg_a = o5_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010110110111",
--  (1139) multiplication_with_reduction_special_prime_3_137
-- reg_a = a6_X; reg_b = b4_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001110000000000100000000000100100010011000011",
--  (1140) multiplication_with_reduction_special_prime_3_138
-- reg_a = o6_X; reg_b = primeSP4; reg_acc = reg_o; o3_X = reg_o; operation : a*b + acc;
"000000100001110000010000100000000000010001110011010111",
--  (1141) multiplication_with_reduction_special_prime_3_139
-- reg_a = a5_X; reg_b = b6_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001110000000000100000100001000100011010100011",
--  (1142) multiplication_with_reduction_special_prime_3_140
-- reg_a = o5_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100011010110111",
--  (1143) multiplication_with_reduction_special_prime_3_141
-- reg_a = a6_X; reg_b = b5_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001110000000000100000000000100100010111000011",
--  (1144) multiplication_with_reduction_special_prime_3_142
-- reg_a = o6_X; reg_b = primeSP5; reg_acc = reg_o; o4_X = reg_o; operation : a*b + acc;
"000000100001110000010000100000000000010110010111010111",
--  (1145) multiplication_with_reduction_special_prime_3_143
-- reg_a = a6_X; reg_b = b6_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001110000000000100000100001100100011011000011",
--  (1146) multiplication_with_reduction_special_prime_3_144
-- reg_a = o6_X; reg_b = primeSP6; reg_acc = reg_o; o5_X = reg_o; o6_X = reg_o >> 256; operation : a*b + acc;
"000000100001110001110000100000000000011010111011010111",
--  (1147) multiplication_with_reduction_special_prime_3_145
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (1148) multiplication_with_reduction_special_prime_3_146
-- -- In case of size 8
-- reg_a = a0_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011000000011",
--  (1149) multiplication_with_reduction_special_prime_3_147
-- reg_a = a6_X; reg_b = b0_X; reg_acc = reg_o; o6_X = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000011111000011000011",
--  (1150) multiplication_with_reduction_special_prime_3_148
-- reg_a = o0_X; reg_b = primeSP7; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001111000000000100000100000000100011100010111",
--  (1151) multiplication_with_reduction_special_prime_3_149
-- reg_a = a1_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011000100011",
--  (1152) multiplication_with_reduction_special_prime_3_150
-- reg_a = o1_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011000110111",
--  (1153) multiplication_with_reduction_special_prime_3_151
-- reg_a = a2_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010101000011",
--  (1154) multiplication_with_reduction_special_prime_3_152
-- reg_a = o2_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010101010111",
--  (1155) multiplication_with_reduction_special_prime_3_153
-- reg_a = a3_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010001100011",
--  (1156) multiplication_with_reduction_special_prime_3_154
-- reg_a = o3_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010001110111",
--  (1157) multiplication_with_reduction_special_prime_3_155
-- reg_a = a4_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001110000011",
--  (1158) multiplication_with_reduction_special_prime_3_156
-- reg_a = o4_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001110010111",
--  (1159) multiplication_with_reduction_special_prime_3_157
-- reg_a = a5_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001010100011",
--  (1160) multiplication_with_reduction_special_prime_3_158
-- reg_a = a6_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100000111000011",
--  (1161) multiplication_with_reduction_special_prime_3_159
-- reg_a = a0_X; reg_b = b7_X; reg_acc = reg_o; Enable sign b; operation : a*b + acc;
"000000100001111000000000100000000001000100011100000011",
--  (1162) multiplication_with_reduction_special_prime_3_160
-- reg_a = a7_X; reg_b = b0_X; reg_acc = reg_o; o7_X = reg_o; Enable sign a; operation : a*b + acc;
"000000100001111000010000100000000000100011100011100011",
--  (1163) multiplication_with_reduction_special_prime_3_161
-- reg_a = a1_X; reg_b = b7_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001111000000000100000100001000100011100100011",
--  (1164) multiplication_with_reduction_special_prime_3_162
-- reg_a = o1_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011100110111",
--  (1165) multiplication_with_reduction_special_prime_3_163
-- reg_a = a2_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011001000011",
--  (1166) multiplication_with_reduction_special_prime_3_164
-- reg_a = o2_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011001010111",
--  (1167) multiplication_with_reduction_special_prime_3_165
-- reg_a = a3_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010101100011",
--  (1168) multiplication_with_reduction_special_prime_3_166
-- reg_a = o3_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010101110111",
--  (1169) multiplication_with_reduction_special_prime_3_167
-- reg_a = a4_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010010000011",
--  (1170) multiplication_with_reduction_special_prime_3_168
-- reg_a = o4_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010010010111",
--  (1171) multiplication_with_reduction_special_prime_3_169
-- reg_a = a5_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001110100011",
--  (1172) multiplication_with_reduction_special_prime_3_170
-- reg_a = o5_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001110110111",
--  (1173) multiplication_with_reduction_special_prime_3_171
-- reg_a = a6_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001011000011",
--  (1174) multiplication_with_reduction_special_prime_3_172
-- reg_a = a7_X; reg_b = b1_X; reg_acc = reg_o; o0_X = reg_o; Enable sign a; operation : a*b + acc;
"000000100001111000010000100000000000100100000111100011",
--  (1175) multiplication_with_reduction_special_prime_3_173
-- reg_a = a2_X; reg_b = b7_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001111000000000100000100001000100011101000011",
--  (1176) multiplication_with_reduction_special_prime_3_174
-- reg_a = o2_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011101010111",
--  (1177) multiplication_with_reduction_special_prime_3_175
-- reg_a = a3_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011001100011",
--  (1178) multiplication_with_reduction_special_prime_3_176
-- reg_a = o3_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011001110111",
--  (1179) multiplication_with_reduction_special_prime_3_177
-- reg_a = a4_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010110000011",
--  (1180) multiplication_with_reduction_special_prime_3_178
-- reg_a = o4_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010110010111",
--  (1181) multiplication_with_reduction_special_prime_3_179
-- reg_a = a5_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010010100011",
--  (1182) multiplication_with_reduction_special_prime_3_180
-- reg_a = o5_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010010110111",
--  (1183) multiplication_with_reduction_special_prime_3_181
-- reg_a = a6_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001111000011",
--  (1184) multiplication_with_reduction_special_prime_3_182
-- reg_a = o6_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001111010111",
--  (1185) multiplication_with_reduction_special_prime_3_183
-- reg_a = a7_X; reg_b = b2_X; reg_acc = reg_o; o1_X = reg_o; Enable sign a; operation : a*b + acc;
"000000100001111000010000100000000000101000101011100011",
--  (1186) multiplication_with_reduction_special_prime_3_184
-- reg_a = a3_X; reg_b = b7_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001111000000000100000100001000100011101100011",
--  (1187) multiplication_with_reduction_special_prime_3_185
-- reg_a = o3_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011101110111",
--  (1188) multiplication_with_reduction_special_prime_3_186
-- reg_a = a4_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011010000011",
--  (1189) multiplication_with_reduction_special_prime_3_187
-- reg_a = o4_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011010010111",
--  (1190) multiplication_with_reduction_special_prime_3_188
-- reg_a = a5_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010110100011",
--  (1191) multiplication_with_reduction_special_prime_3_189
-- reg_a = o5_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010110110111",
--  (1192) multiplication_with_reduction_special_prime_3_190
-- reg_a = a6_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010011000011",
--  (1193) multiplication_with_reduction_special_prime_3_191
-- reg_a = o6_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010011010111",
--  (1194) multiplication_with_reduction_special_prime_3_192
-- reg_a = a7_X; reg_b = b3_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001111000000000100000000000100100001111100011",
--  (1195) multiplication_with_reduction_special_prime_3_193
-- reg_a = o7_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000001101001111110111",
--  (1196) multiplication_with_reduction_special_prime_3_194
-- reg_a = a4_X; reg_b = b7_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001111000000000100000100001000100011110000011",
--  (1197) multiplication_with_reduction_special_prime_3_195
-- reg_a = o4_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011110010111",
--  (1198) multiplication_with_reduction_special_prime_3_196
-- reg_a = a5_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011010100011",
--  (1199) multiplication_with_reduction_special_prime_3_197
-- reg_a = o5_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011010110111",
--  (1200) multiplication_with_reduction_special_prime_3_198
-- reg_a = a6_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010111000011",
--  (1201) multiplication_with_reduction_special_prime_3_199
-- reg_a = o6_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010111010111",
--  (1202) multiplication_with_reduction_special_prime_3_200
-- reg_a = a7_X; reg_b = b4_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001111000000000100000000000100100010011100011",
--  (1203) multiplication_with_reduction_special_prime_3_201
-- reg_a = o7_X; reg_b = primeSP4; reg_acc = reg_o; o3_X = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000010001110011110111",
--  (1204) multiplication_with_reduction_special_prime_3_202
-- reg_a = a5_X; reg_b = b7_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001111000000000100000100001000100011110100011",
--  (1205) multiplication_with_reduction_special_prime_3_203
-- reg_a = o5_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011110110111",
--  (1206) multiplication_with_reduction_special_prime_3_204
-- reg_a = a6_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011011000011",
--  (1207) multiplication_with_reduction_special_prime_3_205
-- reg_a = o6_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011011010111",
--  (1208) multiplication_with_reduction_special_prime_3_206
-- reg_a = a7_X; reg_b = b5_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001111000000000100000000000100100010111100011",
--  (1209) multiplication_with_reduction_special_prime_3_207
-- reg_a = o7_X; reg_b = primeSP5; reg_acc = reg_o; o4_X = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000010110010111110111",
--  (1210) multiplication_with_reduction_special_prime_3_208
-- reg_a = a6_X; reg_b = b7_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001111000000000100000100001000100011111000011",
--  (1211) multiplication_with_reduction_special_prime_3_209
-- reg_a = o6_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011111010111",
--  (1212) multiplication_with_reduction_special_prime_3_210
-- reg_a = a7_X; reg_b = b6_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001111000000000100000000000100100011011100011",
--  (1213) multiplication_with_reduction_special_prime_3_211
-- reg_a = o7_X; reg_b = primeSP6; reg_acc = reg_o; o5_X = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000011010111011110111",
--  (1214) multiplication_with_reduction_special_prime_3_212
-- reg_a = a7_X; reg_b = b7_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001111000000000100000100001100100011111100011",
--  (1215) multiplication_with_reduction_special_prime_3_213
-- reg_a = o7_X; reg_b = primeSP7; reg_acc = reg_o; o6_X = reg_o; o7_X = reg_o >> 256; operation : a*b + acc;
"000000100001111001110000100000000000011111011111110111",
--  (1216) multiplication_with_reduction_special_prime_3_214
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (1217) square_with_reduction_0
-- -- In case of size 1
-- reg_a = a0_X; reg_b = a0_X; reg_acc = 0; Enable sign a,b; operation : a*b + acc;
"000000100001000000000000100000010001100100000000000011",
--  (1218) square_with_reduction_1
-- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o0_X = reg_y; operation : keep accumulator;
"000000100001000000011000110000000100000100000000011011",
--  (1219) square_with_reduction_2
-- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
"000000100001000000000000100000000010000100000000010011",
--  (1220) square_with_reduction_3
-- reg_a = 0; reg_b = 0; reg_acc = reg_o >> 256; o0_X = reg_o; operation : a*b + acc;
"000000100001000000010000100000101110000100000000000011",
--  (1221) square_with_reduction_4
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (1222) square_with_reduction_5
-- -- In case of 2, 3, 4, 5, 6, 7, 8
-- reg_a = a0_X; reg_b = a0_X; reg_acc = 0; operation : a*b + acc;
"000000100001001000000000100000010000000100000000000011",
--  (1223) square_with_reduction_6
-- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o0_X = reg_y; operation : keep accumulator;
"000000100001001000011000110000000100000100000000011011",
--  (1224) square_with_reduction_7
-- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
"000000100001001000000000100000000010000100000000010011",
--  (1225) square_with_reduction_8
-- reg_a = o0_X; reg_b = prime1; reg_acc = reg_o >> 256; operation : a*b + acc;
"000011100001001000000000100000100000000100000100010111",
--  (1226) square_with_reduction_9
-- -- In case of size 2
-- reg_a = a0_X; reg_b = a1_X; reg_acc = reg_o; Enable sign b; operation : 2*a*b + acc;
"000000100001001000000100100000000001000100000100000011",
--  (1227) square_with_reduction_10
-- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o1_X = reg_y; operation : keep accumulator;
"000000100001001000011000110000000100001000100000111011",
--  (1228) square_with_reduction_11
-- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
"000000100001001000000000100000000010000100000000110011",
--  (1229) square_with_reduction_12
-- reg_a = a1_X; reg_b = a1_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001001000000000100000100001100100000100100011",
--  (1230) square_with_reduction_13
-- reg_a = o1_X; reg_b = prime1; reg_acc = reg_o; o0_X = reg_o; o1_X = reg_o >> 256; operation : a*b + acc;
"000000100001001001110000100000000000000100000100110111",
--  (1231) square_with_reduction_14
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (1232) square_with_reduction_15
-- -- Others cases
-- reg_a = a0_X; reg_b = a1_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001010000000100100000000000000100000100000011",
--  (1233) square_with_reduction_16
-- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o1_X = reg_y; operation : keep accumulator;
"000000100001010000011000110000000100001000100000011011",
--  (1234) square_with_reduction_17
-- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
"000000100001010000000000100000000010000100000000010011",
--  (1235) square_with_reduction_18
-- reg_a = o0_X; reg_b = prime2; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001010000000000100000100000000100001000010111",
--  (1236) square_with_reduction_19
-- reg_a = a1_X; reg_b = a1_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001010000000000100000000000000100000100100011",
--  (1237) square_with_reduction_20
-- reg_a = o1_X; reg_b = prime1; reg_acc = reg_o; operation : a*b + acc;
"000101000001010000000000100000000000000100000100110111",
--  (1238) square_with_reduction_21
-- -- In case of size 3
-- reg_a = a0_X; reg_b = a2_X; reg_acc = reg_o; Enable sign b; operation : 2*a*b + acc;
"000000100001010000000100100000000001000100001000000011",
--  (1239) square_with_reduction_22
-- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o2_X = reg_y; operation : keep accumulator;
"000000100001010000011000110000000100001101000000011011",
--  (1240) square_with_reduction_23
-- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
"000000100001010000000000100000000010000100000000010011",
--  (1241) square_with_reduction_24
-- reg_a = a1_X; reg_b = a2_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001010000000100100000100001000100001000100011",
--  (1242) square_with_reduction_25
-- reg_a = o1_X; reg_b = prime2; reg_acc = reg_o; operation : a*b + acc;
"000000100001010000000000100000000000000100001000110111",
--  (1243) square_with_reduction_26
-- reg_a = o2_X; reg_b = prime1; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
"000000100001010000010000100000000000000100000101010111",
--  (1244) square_with_reduction_27
-- reg_a = a2_X; reg_b = a2_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001010000000000100000100001100100001001000011",
--  (1245) square_with_reduction_28
-- reg_a = o2_X; reg_b = prime2; reg_acc = reg_o; o1_X = reg_o; o2_X = reg_o >> 256; operation : a*b + acc;
"000000100001010001110000100000000000001000101001010111",
--  (1246) square_with_reduction_29
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (1247) square_with_reduction_30
-- -- Other cases
-- reg_a = a0_X; reg_b = a2_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001011000000100100000000000000100001000000011",
--  (1248) square_with_reduction_31
-- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o2_X = reg_y; operation : keep accumulator;
"000000100001011000011000110000000100001101000000011011",
--  (1249) square_with_reduction_32
-- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
"000000100001011000000000100000000010000100000000010011",
--  (1250) square_with_reduction_33
-- reg_a = o0_X; reg_b = prime3; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001011000000000100000100000000100001100010111",
--  (1251) square_with_reduction_34
-- reg_a = a1_X; reg_b = a2_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001011000000100100000000000000100001000100011",
--  (1252) square_with_reduction_35
-- reg_a = o1_X; reg_b = prime2; reg_acc = reg_o; operation : a*b + acc;
"000000100001011000000000100000000000000100001000110111",
--  (1253) square_with_reduction_36
-- reg_a = o2_X; reg_b = prime1; reg_acc = reg_o; operation : a*b + acc;
"000111100001011000000000100000000000000100000101010111",
--  (1254) square_with_reduction_37
-- In case of size 4
-- reg_a = a0_X; reg_b = a3_X; reg_acc = reg_o; Enable sign b; operation : 2*a*b + acc;
"000000100001011000000100100000000001000100001100000011",
--  (1255) square_with_reduction_38
-- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o3_X = reg_y; operation : keep accumulator;
"000000100001011000011000110000000100010001100000011011",
--  (1256) square_with_reduction_39
-- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
"000000100001011000000000100000000010000100000000010011",
--  (1257) square_with_reduction_40
-- reg_a = a1_X; reg_b = a3_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001011000000100100000100001000100001100100011",
--  (1258) square_with_reduction_41
-- reg_a = o1_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
"000000100001011000000000100000000000000100001100110111",
--  (1259) square_with_reduction_42
-- reg_a = a2_X; reg_b = a2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001011000000000100000000000000100001001000011",
--  (1260) square_with_reduction_43
-- reg_a = o2_X; reg_b = prime2; reg_acc = reg_o; operation : a*b + acc;
"000000100001011000000000100000000000000100001001010111",
--  (1261) square_with_reduction_44
-- reg_a = o3_X; reg_b = prime1; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
"000000100001011000010000100000000000000100000101110111",
--  (1262) square_with_reduction_45
-- reg_a = a2_X; reg_b = a3_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001011000000100100000100001000100001101000011",
--  (1263) square_with_reduction_46
-- reg_a = o2_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
"000000100001011000000000100000000000000100001101010111",
--  (1264) square_with_reduction_47
-- reg_a = o3_X; reg_b = prime2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
"000000100001011000010000100000000000001000101001110111",
--  (1265) square_with_reduction_48
-- reg_a = a3_X; reg_b = a3_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001011000000000100000100001100100001101100011",
--  (1266) square_with_reduction_49
-- reg_a = o3_X; reg_b = prime3; reg_acc = reg_o; o2_X = reg_o; o3_X = reg_o >> 256; operation : a*b + acc;
"000000100001011001110000100000000000001101001101110111",
--  (1267) square_with_reduction_50
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (1268) square_with_reduction_51
-- -- Other cases
-- reg_a = a0_X; reg_b = a3_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001100000000100100000000000000100001100000011",
--  (1269) square_with_reduction_52
-- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o3_X = reg_y; operation : keep accumulator;
"000000100001100000011000110000000100010001100000011011",
--  (1270) square_with_reduction_53
-- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000010000100000000010011",
--  (1271) square_with_reduction_54
-- reg_a = o0_X; reg_b = prime4; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001100000000000100000100000000100010000010111",
--  (1272) square_with_reduction_55
-- reg_a = a1_X; reg_b = a3_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001100000000100100000000000000100001100100011",
--  (1273) square_with_reduction_56
-- reg_a = o1_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001100110111",
--  (1274) square_with_reduction_57
-- reg_a = a2_X; reg_b = a2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001001000011",
--  (1275) square_with_reduction_58
-- reg_a = o2_X; reg_b = prime2; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001001010111",
--  (1276) square_with_reduction_59
-- reg_a = o3_X; reg_b = prime1; reg_acc = reg_o; operation : a*b + acc;
"001010100001100000000000100000000000000100000101110111",
--  (1277) square_with_reduction_60
-- -- In case of size 5
-- reg_a = a0_X; reg_b = a4_X; reg_acc = reg_o; Enable sign b; operation : 2*a*b + acc;
"000000100001100000000100100000000001000100010000000011",
--  (1278) square_with_reduction_61
-- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o4_X = reg_y; operation : keep accumulator;
"000000100001100000011000110000000100010110000000011011",
--  (1279) square_with_reduction_62
-- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000010000100000000010011",
--  (1280) square_with_reduction_63
-- reg_a = a1_X; reg_b = a4_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001100000000100100000100001000100010000100011",
--  (1281) square_with_reduction_64
-- reg_a = o1_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100010000110111",
--  (1282) square_with_reduction_65
-- reg_a = a2_X; reg_b = a3_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001100000000100100000000000000100001101000011",
--  (1283) square_with_reduction_66
-- reg_a = o2_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001101010111",
--  (1284) square_with_reduction_67
-- reg_a = o3_X; reg_b = prime2; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001001110111",
--  (1285) square_with_reduction_68
-- reg_a = o4_X; reg_b = prime1; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
"000000100001100000010000100000000000000100000110010111",
--  (1286) square_with_reduction_69
-- reg_a = a2_X; reg_b = a4_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001100000000100100000100001000100010001000011",
--  (1287) square_with_reduction_70
-- reg_a = o2_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100010001010111",
--  (1288) square_with_reduction_71
-- reg_a = a3_X; reg_b = a3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001101100011",
--  (1289) square_with_reduction_72
-- reg_a = o3_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001101110111",
--  (1290) square_with_reduction_73
-- reg_a = o4_X; reg_b = prime2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
"000000100001100000010000100000000000001000101010010111",
--  (1291) square_with_reduction_74
-- reg_a = a3_X; reg_b = a4_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001100000000100100000100001000100010001100011",
--  (1292) square_with_reduction_75
-- reg_a = o3_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100010001110111",
--  (1293) square_with_reduction_76
-- reg_a = o4_X; reg_b = prime3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
"000000100001100000010000100000000000001101001110010111",
--  (1294) square_with_reduction_77
-- reg_a = a4_X; reg_b = a4_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001100000000000100000100001100100010010000011",
--  (1295) square_with_reduction_78
-- reg_a = o4_X; reg_b = prime4; reg_acc = reg_o; o3_X = reg_o; o4_X = reg_o >> 256; operation : a*b + acc;
"000000100001100001110000100000000000010001110010010111",
--  (1296) square_with_reduction_79
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (1297) square_with_reduction_80
-- -- Other cases
-- reg_a = a0_X; reg_b = a4_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001101000000100100000000000000100010000000011",
--  (1298) square_with_reduction_81
-- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o4_X = reg_y; operation : keep accumulator;
"000000100001101000011000110000000100010110000000011011",
--  (1299) square_with_reduction_82
-- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000010000100000000010011",
--  (1300) square_with_reduction_83
-- reg_a = o0_X; reg_b = prime5; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001101000000000100000100000000100010100010111",
--  (1301) square_with_reduction_84
-- reg_a = a1_X; reg_b = a4_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001101000000100100000000000000100010000100011",
--  (1302) square_with_reduction_85
-- reg_a = o1_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010000110111",
--  (1303) square_with_reduction_86
-- reg_a = a2_X; reg_b = a3_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001101000000100100000000000000100001101000011",
--  (1304) square_with_reduction_87
-- reg_a = o2_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001101010111",
--  (1305) square_with_reduction_88
-- reg_a = o3_X; reg_b = prime2; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001001110111",
--  (1306) square_with_reduction_89
-- reg_a = o4_X; reg_b = prime1; reg_acc = reg_o; operation : a*b + acc;
"001110100001101000000000100000000000000100000110010111",
--  (1307) square_with_reduction_90
-- -- In case of size 6
-- reg_a = a0_X; reg_b = a5_X; reg_acc = reg_o; Enable sign b; operation : 2*a*b + acc;
"000000100001101000000100100000000001000100010100000011",
--  (1308) square_with_reduction_91
-- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o5_X = reg_y; operation : keep accumulator;
"000000100001101000011000110000000100011010100000011011",
--  (1309) square_with_reduction_92
-- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000010000100000000010011",
--  (1310) square_with_reduction_93
-- reg_a = a1_X; reg_b = a5_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001101000000100100000100001000100010100100011",
--  (1311) square_with_reduction_94
-- reg_a = o1_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010100110111",
--  (1312) square_with_reduction_95
-- reg_a = a2_X; reg_b = a4_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001101000000100100000000000000100010001000011",
--  (1313) square_with_reduction_96
-- reg_a = o2_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010001010111",
--  (1314) square_with_reduction_97
-- reg_a = a3_X; reg_b = a3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001101100011",
--  (1315) square_with_reduction_98
-- reg_a = o3_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001101110111",
--  (1316) square_with_reduction_99
-- reg_a = o4_X; reg_b = prime2; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001010010111",
--  (1317) square_with_reduction_100
-- reg_a = o5_X; reg_b = prime1; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
"000000100001101000010000100000000000000100000110110111",
--  (1318) square_with_reduction_101
-- reg_a = a2_X; reg_b = a5_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001101000000100100000100001000100010101000011",
--  (1319) square_with_reduction_102
-- reg_a = o2_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010101010111",
--  (1320) square_with_reduction_103
-- reg_a = a3_X; reg_b = a4_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001101000000100100000000000000100010001100011",
--  (1321) square_with_reduction_104
-- reg_a = o3_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010001110111",
--  (1322) square_with_reduction_105
-- reg_a = o4_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001110010111",
--  (1323) square_with_reduction_106
-- reg_a = o5_X; reg_b = prime2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
"000000100001101000010000100000000000001000101010110111",
--  (1324) square_with_reduction_107
-- reg_a = a3_X; reg_b = a5_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001101000000100100000100001000100010101100011",
--  (1325) square_with_reduction_108
-- reg_a = o3_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010101110111",
--  (1326) square_with_reduction_109
-- reg_a = a4_X; reg_b = a4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010010000011",
--  (1327) square_with_reduction_110
-- reg_a = o4_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010010010111",
--  (1328) square_with_reduction_111
-- reg_a = o5_X; reg_b = prime3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
"000000100001101000010000100000000000001101001110110111",
--  (1329) square_with_reduction_112
-- reg_a = a4_X; reg_b = a5_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001101000000100100000100001000100010110000011",
--  (1330) square_with_reduction_113
-- reg_a = o4_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010110010111",
--  (1331) square_with_reduction_114
-- reg_a = o5_X; reg_b = prime4; reg_acc = reg_o; o3_X = reg_o; operation : a*b + acc;
"000000100001101000010000100000000000010001110010110111",
--  (1332) square_with_reduction_115
-- reg_a = a5_X; reg_b = a5_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001101000000000100000100001100100010110100011",
--  (1333) square_with_reduction_116
-- reg_a = o5_X; reg_b = prime5; reg_acc = reg_o; o4_X = reg_o; o5_X = reg_o >> 256; operation : a*b + acc;
"000000100001101001110000100000000000010110010110110111",
--  (1334) square_with_reduction_117
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (1335) square_with_reduction_118
-- -- Other cases
-- reg_a = a0_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001110000000100100000000000000100010100000011",
--  (1336) square_with_reduction_119
-- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o5_X = reg_y; operation : keep accumulator;
"000000100001110000011000110000000100010110100000011011",
--  (1337) square_with_reduction_120
-- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000010000100000000010011",
--  (1338) square_with_reduction_121
-- reg_a = o0_X; reg_b = prime6; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001110000000000100000100000000100011000010111",
--  (1339) square_with_reduction_122
-- reg_a = a1_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001110000000100100000000000000100010100100011",
--  (1340) square_with_reduction_123
-- reg_a = o1_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010100110111",
--  (1341) square_with_reduction_124
-- reg_a = a2_X; reg_b = a4_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001110000000100100000000000000100010001000011",
--  (1342) square_with_reduction_125
-- reg_a = o2_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010001010111",
--  (1343) square_with_reduction_126
-- reg_a = a3_X; reg_b = a3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001101100011",
--  (1344) square_with_reduction_127
-- reg_a = o3_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001101110111",
--  (1345) square_with_reduction_128
-- reg_a = o4_X; reg_b = prime2; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001010010111",
--  (1346) square_with_reduction_129
-- reg_a = o5_X; reg_b = prime1; reg_acc = reg_o; operation : a*b + acc;
"010011000001110000000000100000000000000100000110110111",
--  (1347) square_with_reduction_130
-- -- In case of size 7
-- reg_a = a0_X; reg_b = a6_X; reg_acc = reg_o; Enable sign b; operation : 2*a*b + acc;
"000000100001110000000100100000000001000100011000000011",
--  (1348) square_with_reduction_131
-- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o6_X = reg_y; operation : keep accumulator;
"000000100001110000011000110000000100011111000000011011",
--  (1349) square_with_reduction_132
-- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000010000100000000010011",
--  (1350) square_with_reduction_133
-- reg_a = a1_X; reg_b = a6_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001110000000100100000100001000100011000100011",
--  (1351) square_with_reduction_134
-- reg_a = o1_X; reg_b = prime6; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100011000110111",
--  (1352) square_with_reduction_135
-- reg_a = a2_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001110000000100100000000000000100010101000011",
--  (1353) square_with_reduction_136
-- reg_a = o2_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010101010111",
--  (1354) square_with_reduction_137
-- reg_a = a3_X; reg_b = a4_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001110000000100100000000000000100010001100011",
--  (1355) square_with_reduction_138
-- reg_a = o3_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010001110111",
--  (1356) square_with_reduction_139
-- reg_a = o4_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001110010111",
--  (1357) square_with_reduction_140
-- reg_a = o5_X; reg_b = prime2; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001010110111",
--  (1358) square_with_reduction_141
-- reg_a = o6_X; reg_b = prime1; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
"000000100001110000010000100000000000000100000111010111",
--  (1359) square_with_reduction_142
-- reg_a = a2_X; reg_b = a6_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001110000000100100000100001000100011001000011",
--  (1360) square_with_reduction_143
-- reg_a = o2_X; reg_b = prime6; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100011001010111",
--  (1361) square_with_reduction_144
-- reg_a = a3_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001110000000100100000000000000100010101100011",
--  (1362) square_with_reduction_145
-- reg_a = o3_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010101110111",
--  (1363) square_with_reduction_146
-- reg_a = a4_X; reg_b = a4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010010000011",
--  (1364) square_with_reduction_147
-- reg_a = o4_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010010010111",
--  (1365) square_with_reduction_148
-- reg_a = o5_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001110110111",
--  (1366) square_with_reduction_149
-- reg_a = o6_X; reg_b = prime2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
"000000100001110000010000100000000000001000101011010111",
--  (1367) square_with_reduction_150
-- reg_a = a3_X; reg_b = a6_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001110000000100100000100001000100011001100011",
--  (1368) square_with_reduction_151
-- reg_a = o3_X; reg_b = prime6; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100011001110111",
--  (1369) square_with_reduction_152
-- reg_a = a4_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001110000000100100000000000000100010110000011",
--  (1370) square_with_reduction_153
-- reg_a = o4_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010110010111",
--  (1371) square_with_reduction_154
-- reg_a = o5_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010010110111",
--  (1372) square_with_reduction_155
-- reg_a = o6_X; reg_b = prime3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
"000000100001110000010000100000000000001101001111010111",
--  (1373) square_with_reduction_156
-- reg_a = a4_X; reg_b = a6_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001110000000100100000100001000100011010000011",
--  (1374) square_with_reduction_157
-- reg_a = o4_X; reg_b = prime6; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100011010010111",
--  (1375) square_with_reduction_158
-- reg_a = a5_X; reg_b = a5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010110100011",
--  (1376) square_with_reduction_159
-- reg_a = o5_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010110110111",
--  (1377) square_with_reduction_160
-- reg_a = o6_X; reg_b = prime4; reg_acc = reg_o; o3_X = reg_o; operation : a*b + acc;
"000000100001110000010000100000000000010001110011010111",
--  (1378) square_with_reduction_161
-- reg_a = a5_X; reg_b = a6_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001110000000100100000100001000100011010100011",
--  (1379) square_with_reduction_162
-- reg_a = o5_X; reg_b = prime6; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100011010110111",
--  (1380) square_with_reduction_163
-- reg_a = o6_X; reg_b = prime5; reg_acc = reg_o; o4_X = reg_o; operation : a*b + acc;
"000000100001110000010000100000000000010110010111010111",
--  (1381) square_with_reduction_164
-- reg_a = a6_X; reg_b = a6_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001110000000000100000100001100100011011000011",
--  (1382) square_with_reduction_165
-- reg_a = o6_X; reg_b = prime6; reg_acc = reg_o; o5_X = reg_o; o6_X = reg_o >> 256; operation : a*b + acc;
"000000100001110001110000100000000000011010111011010111",
--  (1383) square_with_reduction_166
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (1384) square_with_reduction_167
-- -- In case of size 8
-- reg_a = a0_X; reg_b = a6_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001111000000100100000000000000100011000000011",
--  (1385) square_with_reduction_168
-- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o6_X = reg_y; operation : keep accumulator;
"000000100001111000011000110000000100011111000000011011",
--  (1386) square_with_reduction_169
-- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000010000100000000010011",
--  (1387) square_with_reduction_170
-- reg_a = o0_X; reg_b = prime7; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001111000000000100000100000000100011100010111",
--  (1388) square_with_reduction_171
-- reg_a = a1_X; reg_b = a6_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001111000000100100000000000000100011000100011",
--  (1389) square_with_reduction_172
-- reg_a = o1_X; reg_b = prime6; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011000110111",
--  (1390) square_with_reduction_173
-- reg_a = a2_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001111000000100100000000000000100010101000011",
--  (1391) square_with_reduction_174
-- reg_a = o2_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010101010111",
--  (1392) square_with_reduction_175
-- reg_a = a3_X; reg_b = a4_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001111000000100100000000000000100010001100011",
--  (1393) square_with_reduction_176
-- reg_a = o3_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010001110111",
--  (1394) square_with_reduction_177
-- reg_a = o4_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001010010111",
--  (1395) square_with_reduction_178
-- reg_a = o5_X; reg_b = prime2; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001010110111",
--  (1396) square_with_reduction_179
-- reg_a = o6_X; reg_b = prime1; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100000111010111",
--  (1397) square_with_reduction_180
-- reg_a = a0_X; reg_b = a7_X; reg_acc = reg_o; Enable sign b; operation : 2*a*b + acc;
"000000100001111000000100100000000001000100011100000011",
--  (1398) square_with_reduction_181
-- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o7_X = reg_y; operation : keep accumulator;
"000000100001111000011000110000000100000011100000011011",
--  (1399) square_with_reduction_182
-- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000010000100000000010011",
--  (1400) square_with_reduction_183
-- reg_a = a1_X; reg_b = a7_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001111000000100100000100001000100011100100011",
--  (1401) square_with_reduction_184
-- reg_a = o1_X; reg_b = prime7; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011100110111",
--  (1402) square_with_reduction_185
-- reg_a = a2_X; reg_b = a6_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001111000000100100000000000000100011001000011",
--  (1403) square_with_reduction_186
-- reg_a = o2_X; reg_b = prime6; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011001010111",
--  (1404) square_with_reduction_187
-- reg_a = a3_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001111000000100100000000000000100010101100011",
--  (1405) square_with_reduction_188
-- reg_a = o3_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010101110111",
--  (1406) square_with_reduction_189
-- reg_a = a4_X; reg_b = a4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010010000011",
--  (1407) square_with_reduction_190
-- reg_a = o4_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010010010111",
--  (1408) square_with_reduction_191
-- reg_a = o5_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001110110111",
--  (1409) square_with_reduction_192
-- reg_a = o6_X; reg_b = prime2; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001011010111",
--  (1410) square_with_reduction_193
-- reg_a = o7_X; reg_b = prime1; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000000100000111110111",
--  (1411) square_with_reduction_194
-- reg_a = a2_X; reg_b = a7_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001111000000100100000100001000100011101000011",
--  (1412) square_with_reduction_195
-- reg_a = o2_X; reg_b = prime7; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011101010111",
--  (1413) square_with_reduction_196
-- reg_a = a3_X; reg_b = a6_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001111000000100100000000000000100011001100011",
--  (1414) square_with_reduction_197
-- reg_a = o3_X; reg_b = prime6; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011001110111",
--  (1415) square_with_reduction_198
-- reg_a = a4_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001111000000100100000000000000100010110000011",
--  (1416) square_with_reduction_199
-- reg_a = o4_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010110010111",
--  (1417) square_with_reduction_200
-- reg_a = o5_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010010110111",
--  (1418) square_with_reduction_201
-- reg_a = o6_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001111010111",
--  (1419) square_with_reduction_202
-- reg_a = o7_X; reg_b = prime2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000001000101011110111",
--  (1420) square_with_reduction_203
-- reg_a = a3_X; reg_b = a7_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001111000000100100000100001000100011101100011",
--  (1421) square_with_reduction_204
-- reg_a = o3_X; reg_b = prime7; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011101110111",
--  (1422) square_with_reduction_205
-- reg_a = a4_X; reg_b = a6_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001111000000100100000000000000100011010000011",
--  (1423) square_with_reduction_206
-- reg_a = o4_X; reg_b = prime6; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011010010111",
--  (1424) square_with_reduction_207
-- reg_a = a5_X; reg_b = a5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010110100011",
--  (1425) square_with_reduction_208
-- reg_a = o5_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010110110111",
--  (1426) square_with_reduction_209
-- reg_a = o6_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010011010111",
--  (1427) square_with_reduction_210
-- reg_a = o7_X; reg_b = prime3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000001101001111110111",
--  (1428) square_with_reduction_211
-- reg_a = a4_X; reg_b = a7_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001111000000100100000100001000100011110000011",
--  (1429) square_with_reduction_212
-- reg_a = o4_X; reg_b = prime7; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011110010111",
--  (1430) square_with_reduction_213
-- reg_a = a5_X; reg_b = a6_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001111000000100100000000000000100011010100011",
--  (1431) square_with_reduction_214
-- reg_a = o5_X; reg_b = prime6; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011010110111",
--  (1432) square_with_reduction_215
-- reg_a = o6_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010111010111",
--  (1433) square_with_reduction_216
-- reg_a = o7_X; reg_b = prime4; reg_acc = reg_o; o3_X = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000010001110011110111",
--  (1434) square_with_reduction_217
-- reg_a = a5_X; reg_b = a7_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001111000000100100000100001000100011110100011",
--  (1435) square_with_reduction_218
-- reg_a = o5_X; reg_b = prime7; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011110110111",
--  (1436) square_with_reduction_219
-- reg_a = a6_X; reg_b = a6_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011011000011",
--  (1437) square_with_reduction_220
-- reg_a = o6_X; reg_b = prime6; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011011010111",
--  (1438) square_with_reduction_221
-- reg_a = o7_X; reg_b = prime5; reg_acc = reg_o; o4_X = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000010110010111110111",
--  (1439) square_with_reduction_222
-- reg_a = a6_X; reg_b = a7_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001111000000100100000100001000100011111000011",
--  (1440) square_with_reduction_223
-- reg_a = o6_X; reg_b = prime7; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011111010111",
--  (1441) square_with_reduction_224
-- reg_a = o7_X; reg_b = prime6; reg_acc = reg_o; o5_X = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000011010111011110111",
--  (1442) square_with_reduction_225
-- reg_a = a7_X; reg_b = a7_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001111000000000100000100001100100011111100011",
--  (1443) square_with_reduction_226
-- reg_a = o7_X; reg_b = prime7; reg_acc = reg_o; o6_X = reg_o; o7_X = reg_o >> 256; operation : a*b + acc;
"000000100001111001110000100000000000011111011111110111",
--  (1444) square_with_reduction_227
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (1445) square_with_reduction_special_prime_1_0
-- -- In case of size 1
-- reg_a = a0_X; reg_b = a0_X; reg_acc = 0; Enable sign a,b; operation : a*b + acc;
"000000100001000000000000100000010001100100000000000011",
--  (1446) square_with_reduction_special_prime_1_1
-- reg_a = 0; reg_b = 0; reg_acc = reg_o >> 256; o0_X = reg_o; operation : a*b + acc;
"000000100001000000010000100000101110000100000000000011",
--  (1447) square_with_reduction_special_prime_1_2
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (1448) square_with_reduction_special_prime_1_3
-- -- In case of size 2, 3, 4, 5, 6, 7, 8
-- reg_a = a0_X; reg_b = a0_X; reg_acc = 0; o0_X = reg_o; operation : a*b + acc;
"000000100001001000010000100000010000000100000000000011",
--  (1449) square_with_reduction_special_prime_1_4
-- reg_a = reg_o; reg_b = primeSP1; reg_acc = reg_o >> 256; operation : a*b + acc;
"000010100001001000000000100000100100001000100100010111",
--  (1450) square_with_reduction_special_prime_1_5
-- -- In case of size 2
-- reg_a = a0_X; reg_b = a1_X; reg_acc = reg_o; o1_X = reg_o; Enable sign b; operation : 2*a*b + acc;
"000000100001001000010100100000000001001000100100000011",
--  (1451) square_with_reduction_special_prime_1_6
-- reg_a = a1_X; reg_b = a1_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001001000000000100000100001100100000100100011",
--  (1452) square_with_reduction_special_prime_1_7
-- reg_a = o1_X; reg_b = primeSP1; reg_acc = reg_o; o0_X = reg_o; o1_X = reg_o >> 256; operation : a*b + acc;
"000000100001001001110000100000000000000100000100110111",
--  (1453) square_with_reduction_special_prime_1_8
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (1454) square_with_reduction_special_prime_1_9
-- -- In case of size 3, 4, 5, 6, 7, 8
-- reg_a = a0_X; reg_b = a1_X; reg_acc = reg_o; o1_X = reg_o; operation : 2*a*b + acc;
"000000100001010000010100100000000000001000100100000011",
--  (1455) square_with_reduction_special_prime_1_10
-- reg_a = o0_X; reg_b = primeSP2; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001010000000000100000100000000100001000010111",
--  (1456) square_with_reduction_special_prime_1_11
-- reg_a = a1_X; reg_b = a1_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001010000000000100000000000000100000100100011",
--  (1457) square_with_reduction_special_prime_1_12
-- reg_a = o1_X; reg_b = primeSP1; reg_acc = reg_o; operation : a*b + acc;
"000100000001010000000000100000000000001101000100110111",
--  (1458) square_with_reduction_special_prime_1_13
-- -- In case of size 3
-- reg_a = a0_X; reg_b = a2_X; reg_acc = reg_o; o2_X = reg_o; Enable sign b; operation : 2*a*b + acc;
"000000100001010000010100100000000001001101001000000011",
--  (1459) square_with_reduction_special_prime_1_14
-- reg_a = a1_X; reg_b = a2_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001010000000100100000100001000100001000100011",
--  (1460) square_with_reduction_special_prime_1_15
-- reg_a = o1_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
"000000100001010000000000100000000000000100001000110111",
--  (1461) square_with_reduction_special_prime_1_16
-- reg_a = o2_X; reg_b = primeSP1; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
"000000100001010000010000100000000000000100000101010111",
--  (1462) square_with_reduction_special_prime_1_17
-- reg_a = a2_X; reg_b = a2_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001010000000000100000100001100100001001000011",
--  (1463) square_with_reduction_special_prime_1_18
-- reg_a = o2_X; reg_b = primeSP2; reg_acc = reg_o; o1_X = reg_o; o2_X = reg_o >> 256; operation : a*b + acc;
"000000100001010001110000100000000000001000101001010111",
--  (1464) square_with_reduction_special_prime_1_19
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (1465) square_with_reduction_special_prime_1_20
-- -- In case of sizes 4, 5, 6, 7, 8
-- reg_a = a0_X; reg_b = a2_X; reg_acc = reg_o; o2_X = reg_o; operation : 2*a*b + acc;
"000000100001011000010100100000000000001101001000000011",
--  (1466) square_with_reduction_special_prime_1_21
-- reg_a = o0_X; reg_b = primeSP3; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001011000000000100000100000000100001100010111",
--  (1467) square_with_reduction_special_prime_1_22
-- reg_a = a1_X; reg_b = a2_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001011000000100100000000000000100001000100011",
--  (1468) square_with_reduction_special_prime_1_23
-- reg_a = o1_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
"000000100001011000000000100000000000000100001000110111",
--  (1469) square_with_reduction_special_prime_1_24
-- reg_a = o2_X; reg_b = primeSP1; reg_acc = reg_o; operation : a*b + acc;
"000110100001011000000000100000000000000100000101010111",
--  (1470) square_with_reduction_special_prime_1_25
-- -- In case of size 4
-- reg_a = a0_X; reg_b = a3_X; reg_acc = reg_o; o3_X = reg_o; Enable sign b; operation : 2*a*b + acc;
"000000100001011000010100100000000001010001101100000011",
--  (1471) square_with_reduction_special_prime_1_26
-- reg_a = a1_X; reg_b = a3_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001011000000100100000100001000100001100100011",
--  (1472) square_with_reduction_special_prime_1_27
-- reg_a = o1_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001011000000000100000000000000100001100110111",
--  (1473) square_with_reduction_special_prime_1_28
-- reg_a = a2_X; reg_b = a2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001011000000000100000000000000100001001000011",
--  (1474) square_with_reduction_special_prime_1_29
-- reg_a = o2_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
"000000100001011000000000100000000000000100001001010111",
--  (1475) square_with_reduction_special_prime_1_30
-- reg_a = o3_X; reg_b = primeSP1; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
"000000100001011000010000100000000000000100000101110111",
--  (1476) square_with_reduction_special_prime_1_31
-- reg_a = a2_X; reg_b = a3_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001011000000100100000100001000100001101000011",
--  (1477) square_with_reduction_special_prime_1_32
-- reg_a = o2_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001011000000000100000000000000100001101010111",
--  (1478) square_with_reduction_special_prime_1_33
-- reg_a = o3_X; reg_b = primeSP2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
"000000100001011000010000100000000000001000101001110111",
--  (1479) square_with_reduction_special_prime_1_34
-- reg_a = a3_X; reg_b = a3_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001011000000000100000100001100100001101100011",
--  (1480) square_with_reduction_special_prime_1_35
-- reg_a = o3_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; o3_X = reg_o >> 256; operation : a*b + acc;
"000000100001011001110000100000000000001101001101110111",
--  (1481) square_with_reduction_special_prime_1_36
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (1482) square_with_reduction_special_prime_1_37
-- -- In case of sizes 5, 6, 7, 8
-- reg_a = a0_X; reg_b = a3_X; reg_acc = reg_o; o3_X = reg_o; operation : 2*a*b + acc;
"000000100001100000010100100000000000010001101100000011",
--  (1483) square_with_reduction_special_prime_1_38
-- reg_a = o0_X; reg_b = primeSP4; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001100000000000100000100000000100010000010111",
--  (1484) square_with_reduction_special_prime_1_39
-- reg_a = a1_X; reg_b = a3_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001100000000100100000000000000100001100100011",
--  (1485) square_with_reduction_special_prime_1_40
-- reg_a = o1_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001100110111",
--  (1486) square_with_reduction_special_prime_1_41
-- reg_a = a2_X; reg_b = a2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001001000011",
--  (1487) square_with_reduction_special_prime_1_42
-- reg_a = o2_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001001010111",
--  (1488) square_with_reduction_special_prime_1_43
-- reg_a = o3_X; reg_b = primeSP1; reg_acc = reg_o; operation : a*b + acc;
"001001100001100000000000100000000000000100000101110111",
--  (1489) square_with_reduction_special_prime_1_44
-- -- In case of size 5
-- reg_a = a0_X; reg_b = a4_X; reg_acc = reg_o; o4_X = reg_o; Enable sign b; operation : 2*a*b + acc;
"000000100001100000010100100000000001010110010000000011",
--  (1490) square_with_reduction_special_prime_1_45
-- reg_a = a1_X; reg_b = a4_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001100000000100100000100001000100010000100011",
--  (1491) square_with_reduction_special_prime_1_46
-- reg_a = o1_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100010000110111",
--  (1492) square_with_reduction_special_prime_1_47
-- reg_a = a2_X; reg_b = a3_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001100000000100100000000000000100001101000011",
--  (1493) square_with_reduction_special_prime_1_48
-- reg_a = o2_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001101010111",
--  (1494) square_with_reduction_special_prime_1_49
-- reg_a = o3_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001001110111",
--  (1495) square_with_reduction_special_prime_1_50
-- reg_a = o4_X; reg_b = primeSP1; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
"000000100001100000010000100000000000000100000110010111",
--  (1496) square_with_reduction_special_prime_1_51
-- reg_a = a2_X; reg_b = a4_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001100000000100100000100001000100010001000011",
--  (1497) square_with_reduction_special_prime_1_52
-- reg_a = o2_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100010001010111",
--  (1498) square_with_reduction_special_prime_1_53
-- reg_a = a3_X; reg_b = a3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001101100011",
--  (1499) square_with_reduction_special_prime_1_54
-- reg_a = o3_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001101110111",
--  (1500) square_with_reduction_special_prime_1_55
-- reg_a = o4_X; reg_b = primeSP2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
"000000100001100000010000100000000000001000101010010111",
--  (1501) square_with_reduction_special_prime_1_56
-- reg_a = a3_X; reg_b = a4_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001100000000100100000100001000100010001100011",
--  (1502) square_with_reduction_special_prime_1_57
-- reg_a = o3_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100010001110111",
--  (1503) square_with_reduction_special_prime_1_58
-- reg_a = o4_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
"000000100001100000010000100000000000001101001110010111",
--  (1504) square_with_reduction_special_prime_1_59
-- reg_a = a4_X; reg_b = a4_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001100000000000100000100001100100010010000011",
--  (1505) square_with_reduction_special_prime_1_60
-- reg_a = o4_X; reg_b = primeSP4; reg_acc = reg_o; o3_X = reg_o; o4_X = reg_o >> 256; operation : a*b + acc;
"000000100001100001110000100000000000010001110010010111",
--  (1506) square_with_reduction_special_prime_1_61
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (1507) square_with_reduction_special_prime_1_62
-- -- In case of sizes 6, 7, 8
-- reg_a = a0_X; reg_b = a4_X; reg_acc = reg_o; o4_X = reg_o; operation : 2*a*b + acc;
"000000100001101000010100100000000000010110010000000011",
--  (1508) square_with_reduction_special_prime_1_63
-- reg_a = o0_X; reg_b = primeSP5; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001101000000000100000100000000100010100010111",
--  (1509) square_with_reduction_special_prime_1_64
-- reg_a = a1_X; reg_b = a4_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001101000000100100000000000000100010000100011",
--  (1510) square_with_reduction_special_prime_1_65
-- reg_a = o1_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010000110111",
--  (1511) square_with_reduction_special_prime_1_66
-- reg_a = a2_X; reg_b = a3_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001101000000100100000000000000100001101000011",
--  (1512) square_with_reduction_special_prime_1_67
-- reg_a = o2_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001101010111",
--  (1513) square_with_reduction_special_prime_1_68
-- reg_a = o3_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001001110111",
--  (1514) square_with_reduction_special_prime_1_69
-- reg_a = o4_X; reg_b = primeSP1; reg_acc = reg_o; operation : a*b + acc;
"001101100001101000000000100000000000000100000110010111",
--  (1515) square_with_reduction_special_prime_1_70
-- -- In case of size 6
-- reg_a = a0_X; reg_b = a5_X; reg_acc = reg_o; o5_X = reg_o; Enable sign b; operation : 2*a*b + acc;
"000000100001101000010100100000000001010010110100000011",
--  (1516) square_with_reduction_special_prime_1_71
-- reg_a = a1_X; reg_b = a5_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001101000000100100000100001000100010100100011",
--  (1517) square_with_reduction_special_prime_1_72
-- reg_a = o1_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010100110111",
--  (1518) square_with_reduction_special_prime_1_73
-- reg_a = a2_X; reg_b = a4_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001101000000100100000000000000100010001000011",
--  (1519) square_with_reduction_special_prime_1_74
-- reg_a = o2_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010001010111",
--  (1520) square_with_reduction_special_prime_1_75
-- reg_a = a3_X; reg_b = a3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001101100011",
--  (1521) square_with_reduction_special_prime_1_76
-- reg_a = o3_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001101110111",
--  (1522) square_with_reduction_special_prime_1_77
-- reg_a = o4_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001010010111",
--  (1523) square_with_reduction_special_prime_1_78
-- reg_a = o5_X; reg_b = primeSP1; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
"000000100001101000010000100000000000000100000110110111",
--  (1524) square_with_reduction_special_prime_1_79
-- reg_a = a2_X; reg_b = a5_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001101000000100100000100001000100010101000011",
--  (1525) square_with_reduction_special_prime_1_80
-- reg_a = o2_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010101010111",
--  (1526) square_with_reduction_special_prime_1_81
-- reg_a = a3_X; reg_b = a4_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001101000000100100000000000000100010001100011",
--  (1527) square_with_reduction_special_prime_1_82
-- reg_a = o3_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010001110111",
--  (1528) square_with_reduction_special_prime_1_83
-- reg_a = o4_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001110010111",
--  (1529) square_with_reduction_special_prime_1_84
-- reg_a = o5_X; reg_b = primeSP2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
"000000100001101000010000100000000000001000101010110111",
--  (1530) square_with_reduction_special_prime_1_85
-- reg_a = a3_X; reg_b = a5_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001101000000100100000100001000100010101100011",
--  (1531) square_with_reduction_special_prime_1_86
-- reg_a = o3_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010101110111",
--  (1532) square_with_reduction_special_prime_1_87
-- reg_a = a4_X; reg_b = a4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010010000011",
--  (1533) square_with_reduction_special_prime_1_88
-- reg_a = o4_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010010010111",
--  (1534) square_with_reduction_special_prime_1_89
-- reg_a = o5_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
"000000100001101000010000100000000000001101001110110111",
--  (1535) square_with_reduction_special_prime_1_90
-- reg_a = a4_X; reg_b = a5_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001101000000100100000100001000100010110000011",
--  (1536) square_with_reduction_special_prime_1_91
-- reg_a = o4_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010110010111",
--  (1537) square_with_reduction_special_prime_1_92
-- reg_a = o5_X; reg_b = primeSP4; reg_acc = reg_o; o3_X = reg_o; operation : a*b + acc;
"000000100001101000010000100000000000010001110010110111",
--  (1538) square_with_reduction_special_prime_1_93
-- reg_a = a5_X; reg_b = a5_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001101000000000100000100001100100010110100011",
--  (1539) square_with_reduction_special_prime_1_94
-- reg_a = o5_X; reg_b = primeSP5; reg_acc = reg_o; o4_X = reg_o; o5_X = reg_o >> 256; operation : a*b + acc;
"000000100001101001110000100000000000010110010110110111",
--  (1540) square_with_reduction_special_prime_1_95
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (1541) square_with_reduction_special_prime_1_96
-- -- In case of sizes 7, 8
-- reg_a = a0_X; reg_b = a5_X; reg_acc = reg_o; o5_X = reg_o; operation : 2*a*b + acc;
"000000100001110000010100100000000000011010110100000011",
--  (1542) square_with_reduction_special_prime_1_97
-- reg_a = o0_X; reg_b = primeSP6; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001110000000000100000100000000100011000010111",
--  (1543) square_with_reduction_special_prime_1_98
-- reg_a = a1_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001110000000100100000000000000100010100100011",
--  (1544) square_with_reduction_special_prime_1_99
-- reg_a = o1_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010100110111",
--  (1545) square_with_reduction_special_prime_1_100
-- reg_a = a2_X; reg_b = a4_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001110000000100100000000000000100010001000011",
--  (1546) square_with_reduction_special_prime_1_101
-- reg_a = o2_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010001010111",
--  (1547) square_with_reduction_special_prime_1_102
-- reg_a = a3_X; reg_b = a3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001101100011",
--  (1548) square_with_reduction_special_prime_1_103
-- reg_a = o3_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001101110111",
--  (1549) square_with_reduction_special_prime_1_104
-- reg_a = o4_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001010010111",
--  (1550) square_with_reduction_special_prime_1_105
-- reg_a = o5_X; reg_b = primeSP1; reg_acc = reg_o; operation : a*b + acc;
"010010000001110000000000100000000000000100000110110111",
--  (1551) square_with_reduction_special_prime_1_106
-- -- In case of size 7
-- reg_a = a0_X; reg_b = a6_X; reg_acc = reg_o; o6_X = reg_o; Enable sign b; operation : 2*a*b + acc;
"000000100001110000010100100000000001011111011000000011",
--  (1552) square_with_reduction_special_prime_1_107
-- reg_a = a1_X; reg_b = a6_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001110000000100100000100001000100011000100011",
--  (1553) square_with_reduction_special_prime_1_108
-- reg_a = o1_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100011000110111",
--  (1554) square_with_reduction_special_prime_1_109
-- reg_a = a2_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001110000000100100000000000000100010101000011",
--  (1555) square_with_reduction_special_prime_1_110
-- reg_a = o2_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010101010111",
--  (1556) square_with_reduction_special_prime_1_111
-- reg_a = a3_X; reg_b = a4_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001110000000100100000000000000100010001100011",
--  (1557) square_with_reduction_special_prime_1_112
-- reg_a = o3_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010001110111",
--  (1558) square_with_reduction_special_prime_1_113
-- reg_a = o4_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001110010111",
--  (1559) square_with_reduction_special_prime_1_114
-- reg_a = o5_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001010110111",
--  (1560) square_with_reduction_special_prime_1_115
-- reg_a = o6_X; reg_b = primeSP1; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
"000000100001110000010000100000000000000100000111010111",
--  (1561) square_with_reduction_special_prime_1_116
-- reg_a = a2_X; reg_b = a6_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001110000000100100000100001000100011001000011",
--  (1562) square_with_reduction_special_prime_1_117
-- reg_a = o2_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100011001010111",
--  (1563) square_with_reduction_special_prime_1_118
-- reg_a = a3_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001110000000100100000000000000100010101100011",
--  (1564) square_with_reduction_special_prime_1_119
-- reg_a = o3_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010101110111",
--  (1565) square_with_reduction_special_prime_1_120
-- reg_a = a4_X; reg_b = a4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010010000011",
--  (1566) square_with_reduction_special_prime_1_121
-- reg_a = o4_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010010010111",
--  (1567) square_with_reduction_special_prime_1_122
-- reg_a = o5_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001110110111",
--  (1568) square_with_reduction_special_prime_1_123
-- reg_a = o6_X; reg_b = primeSP2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
"000000100001110000010000100000000000001000101011010111",
--  (1569) square_with_reduction_special_prime_1_124
-- reg_a = a3_X; reg_b = a6_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001110000000100100000100001000100011001100011",
--  (1570) square_with_reduction_special_prime_1_125
-- reg_a = o3_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100011001110111",
--  (1571) square_with_reduction_special_prime_1_126
-- reg_a = a4_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001110000000100100000000000000100010110000011",
--  (1572) square_with_reduction_special_prime_1_127
-- reg_a = o4_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010110010111",
--  (1573) square_with_reduction_special_prime_1_128
-- reg_a = o5_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010010110111",
--  (1574) square_with_reduction_special_prime_1_129
-- reg_a = o6_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
"000000100001110000010000100000000000001101001111010111",
--  (1575) square_with_reduction_special_prime_1_130
-- reg_a = a4_X; reg_b = a6_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001110000000100100000100001000100011010000011",
--  (1576) square_with_reduction_special_prime_1_131
-- reg_a = o4_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100011010010111",
--  (1577) square_with_reduction_special_prime_1_132
-- reg_a = a5_X; reg_b = a5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010110100011",
--  (1578) square_with_reduction_special_prime_1_133
-- reg_a = o5_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010110110111",
--  (1579) square_with_reduction_special_prime_1_134
-- reg_a = o6_X; reg_b = primeSP4; reg_acc = reg_o; o3_X = reg_o; operation : a*b + acc;
"000000100001110000010000100000000000010001110011010111",
--  (1580) square_with_reduction_special_prime_1_135
-- reg_a = a5_X; reg_b = a6_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001110000000100100000100001000100011010100011",
--  (1581) square_with_reduction_special_prime_1_136
-- reg_a = o5_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100011010110111",
--  (1582) square_with_reduction_special_prime_1_137
-- reg_a = o6_X; reg_b = primeSP5; reg_acc = reg_o; o4_X = reg_o; operation : a*b + acc;
"000000100001110000010000100000000000010110010111010111",
--  (1583) square_with_reduction_special_prime_1_138
-- reg_a = a6_X; reg_b = a6_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001110000000000100000100001100100011011000011",
--  (1584) square_with_reduction_special_prime_1_139
-- reg_a = o6_X; reg_b = primeSP6; reg_acc = reg_o; o5_X = reg_o; o6_X = reg_o >> 256; operation : a*b + acc;
"000000100001110001110000100000000000011010111011010111",
--  (1585) square_with_reduction_special_prime_1_140
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (1586) square_with_reduction_special_prime_1_141
-- -- In case of size 8
-- reg_a = a0_X; reg_b = a6_X; reg_acc = reg_o; o6_X = reg_o; operation : 2*a*b + acc;
"000000100001111000010100100000000000011111011000000011",
--  (1587) square_with_reduction_special_prime_1_142
-- reg_a = o0_X; reg_b = primeSP7; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001111000000000100000100000000100011100010111",
--  (1588) square_with_reduction_special_prime_1_143
-- reg_a = a1_X; reg_b = a6_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001111000000100100000000000000100011000100011",
--  (1589) square_with_reduction_special_prime_1_144
-- reg_a = o1_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011000110111",
--  (1590) square_with_reduction_special_prime_1_145
-- reg_a = a2_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001111000000100100000000000000100010101000011",
--  (1591) square_with_reduction_special_prime_1_146
-- reg_a = o2_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010101010111",
--  (1592) square_with_reduction_special_prime_1_147
-- reg_a = a3_X; reg_b = a4_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001111000000100100000000000000100010001100011",
--  (1593) square_with_reduction_special_prime_1_148
-- reg_a = o3_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010001110111",
--  (1594) square_with_reduction_special_prime_1_149
-- reg_a = o4_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001110010111",
--  (1595) square_with_reduction_special_prime_1_150
-- reg_a = o5_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001010110111",
--  (1596) square_with_reduction_special_prime_1_151
-- reg_a = o6_X; reg_b = primeSP1; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100000111010111",
--  (1597) square_with_reduction_special_prime_1_152
-- reg_a = a0_X; reg_b = a7_X; reg_acc = reg_o; o7_X = reg_o; Enable sign b; operation : 2*a*b + acc;
"000000100001111000010100100000000001000011111100000011",
--  (1598) square_with_reduction_special_prime_1_153
-- reg_a = a1_X; reg_b = a7_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001111000000100100000100001000100011100100011",
--  (1599) square_with_reduction_special_prime_1_154
-- reg_a = o1_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011100110111",
--  (1600) square_with_reduction_special_prime_1_155
-- reg_a = a2_X; reg_b = a6_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001111000000100100000000000000100011001000011",
--  (1601) square_with_reduction_special_prime_1_156
-- reg_a = o2_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011001010111",
--  (1602) square_with_reduction_special_prime_1_157
-- reg_a = a3_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001111000000100100000000000000100010101100011",
--  (1603) square_with_reduction_special_prime_1_158
-- reg_a = o3_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010101110111",
--  (1604) square_with_reduction_special_prime_1_159
-- reg_a = a4_X; reg_b = a4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010010000011",
--  (1605) square_with_reduction_special_prime_1_160
-- reg_a = o4_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010010010111",
--  (1606) square_with_reduction_special_prime_1_161
-- reg_a = o5_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001110110111",
--  (1607) square_with_reduction_special_prime_1_162
-- reg_a = o6_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001011010111",
--  (1608) square_with_reduction_special_prime_1_163
-- reg_a = o7_X; reg_b = primeSP1; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000000100000111110111",
--  (1609) square_with_reduction_special_prime_1_164
-- reg_a = a2_X; reg_b = a7_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001111000000100100000100001000100011101000011",
--  (1610) square_with_reduction_special_prime_1_165
-- reg_a = o2_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011101010111",
--  (1611) square_with_reduction_special_prime_1_166
-- reg_a = a3_X; reg_b = a6_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001111000000100100000000000000100011001100011",
--  (1612) square_with_reduction_special_prime_1_167
-- reg_a = o3_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011001110111",
--  (1613) square_with_reduction_special_prime_1_168
-- reg_a = a4_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001111000000100100000000000000100010110000011",
--  (1614) square_with_reduction_special_prime_1_169
-- reg_a = o4_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010110010111",
--  (1615) square_with_reduction_special_prime_1_170
-- reg_a = o5_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010010110111",
--  (1616) square_with_reduction_special_prime_1_171
-- reg_a = o6_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001111010111",
--  (1617) square_with_reduction_special_prime_1_172
-- reg_a = o7_X; reg_b = primeSP2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000001000101011110111",
--  (1618) square_with_reduction_special_prime_1_173
-- reg_a = a3_X; reg_b = a7_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001111000000100100000100001000100011101100011",
--  (1619) square_with_reduction_special_prime_1_174
-- reg_a = o3_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011101110111",
--  (1620) square_with_reduction_special_prime_1_175
-- reg_a = a4_X; reg_b = a6_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001111000000100100000000000000100011010000011",
--  (1621) square_with_reduction_special_prime_1_176
-- reg_a = o4_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011010010111",
--  (1622) square_with_reduction_special_prime_1_177
-- reg_a = a5_X; reg_b = a5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010110100011",
--  (1623) square_with_reduction_special_prime_1_178
-- reg_a = o5_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010110110111",
--  (1624) square_with_reduction_special_prime_1_179
-- reg_a = o6_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010011010111",
--  (1625) square_with_reduction_special_prime_1_180
-- reg_a = o7_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000001101001111110111",
--  (1626) square_with_reduction_special_prime_1_181
-- reg_a = a4_X; reg_b = a7_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001111000000100100000100001000100011110000011",
--  (1627) square_with_reduction_special_prime_1_182
-- reg_a = o4_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011110010111",
--  (1628) square_with_reduction_special_prime_1_183
-- reg_a = a5_X; reg_b = a6_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001111000000100100000000000000100011010100011",
--  (1629) square_with_reduction_special_prime_1_184
-- reg_a = o5_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011010110111",
--  (1630) square_with_reduction_special_prime_1_185
-- reg_a = o6_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010111010111",
--  (1631) square_with_reduction_special_prime_1_186
-- reg_a = o7_X; reg_b = primeSP4; reg_acc = reg_o; o3_X = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000010001110011110111",
--  (1632) square_with_reduction_special_prime_1_187
-- reg_a = a5_X; reg_b = a7_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001111000000100100000100001000100011110100011",
--  (1633) square_with_reduction_special_prime_1_188
-- reg_a = o5_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011110110111",
--  (1634) square_with_reduction_special_prime_1_189
-- reg_a = a6_X; reg_b = a6_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011011000011",
--  (1635) square_with_reduction_special_prime_1_190
-- reg_a = o6_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011011010111",
--  (1636) square_with_reduction_special_prime_1_191
-- reg_a = o7_X; reg_b = primeSP5; reg_acc = reg_o; o4_X = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000010110010111110111",
--  (1637) square_with_reduction_special_prime_1_192
-- reg_a = a6_X; reg_b = a7_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001111000000100100000100001000100011111000011",
--  (1638) square_with_reduction_special_prime_1_193
-- reg_a = o6_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011111010111",
--  (1639) square_with_reduction_special_prime_1_194
-- reg_a = o7_X; reg_b = primeSP6; reg_acc = reg_o; o5_X = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000011010111011110111",
--  (1640) square_with_reduction_special_prime_1_195
-- reg_a = a7_X; reg_b = a7_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001111000000000100000100001100100011111100011",
--  (1641) square_with_reduction_special_prime_1_196
-- reg_a = o7_X; reg_b = primeSP7; reg_acc = reg_o; o6_X = reg_o; o7_X = reg_o >> 256; operation : a*b + acc;
"000000100001111001110000100000000000011111011111110111",
--  (1642) square_with_reduction_special_prime_1_197
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (1643) square_with_reduction_special_prime_2_0
-- -- In case of size 2, 3, 4, 5, 6, 7, 8
-- reg_a = a0_X; reg_b = a0_X; reg_acc = 0; o0_X = reg_o; operation : a*b + acc;
"000010000001001000010000100000010000000100000000000011",
--  (1644) square_with_reduction_special_prime_2_1
-- -- In case of size 2
-- reg_a = a0_X; reg_b = a1_X; reg_acc = reg_o; o1_X = reg_o; Enable sign b; operation : 2*a*b + acc;
"000000100001001000010100100000000001001000100100000011",
--  (1645) square_with_reduction_special_prime_2_2
-- reg_a = a1_X; reg_b = a1_X; reg_acc = reg_o >> 256; Enable sign a,b; o0_X = reg_o; o1_X = reg_o >> 256; operation : a*b + acc;
"000000100001001001110000100000100001100100000100100011",
--  (1646) square_with_reduction_special_prime_2_3
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (1647) square_with_reduction_special_prime_2_4
-- -- In case of size 3, 4, 5, 6, 7, 8
-- reg_a = a0_X; reg_b = a1_X; reg_acc = reg_o >> 256; o1_X = reg_o; operation : 2*a*b + acc;
"000000100001010000010100100000100000001000100100000011",
--  (1648) square_with_reduction_special_prime_2_5
-- reg_a = o0_X; reg_b = primeSP2; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001010000000000100000100000000100001000010111",
--  (1649) square_with_reduction_special_prime_2_6
-- reg_a = a1_X; reg_b = a1_X; reg_acc = reg_o; operation : a*b + acc;
"000011100001010000000000100000000000000100000100100011",
--  (1650) square_with_reduction_special_prime_2_7
-- -- In case of size 3
-- reg_a = a0_X; reg_b = a2_X; reg_acc = reg_o; o2_X = reg_o; Enable sign b; operation : 2*a*b + acc;
"000000100001010000010100100000000001001101001000000011",
--  (1651) square_with_reduction_special_prime_2_8
-- reg_a = a1_X; reg_b = a2_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001010000000100100000100001000100001000100011",
--  (1652) square_with_reduction_special_prime_2_9
-- reg_a = o1_X; reg_b = primeSP2; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
"000000100001010000010000100000000000000100001000110111",
--  (1653) square_with_reduction_special_prime_2_10
-- reg_a = a2_X; reg_b = a2_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001010000000000100000100001100100001001000011",
--  (1654) square_with_reduction_special_prime_2_11
-- reg_a = o2_X; reg_b = primeSP2; reg_acc = reg_o; o1_X = reg_o; o2_X = reg_o >> 256; operation : a*b + acc;
"000000100001010001110000100000000000001000101001010111",
--  (1655) square_with_reduction_special_prime_2_12
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (1656) square_with_reduction_special_prime_2_13
-- -- In case of size 4, 5, 6, 7, 8
-- reg_a = a0_X; reg_b = a2_X; reg_acc = reg_o; o2_X = reg_o; operation : 2*a*b + acc;
"000000100001011000010100100000000000001101001000000011",
--  (1657) square_with_reduction_special_prime_2_14
-- reg_a = o0_X; reg_b = primeSP3; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001011000000000100000100000000100001100010111",
--  (1658) square_with_reduction_special_prime_2_15
-- reg_a = a1_X; reg_b = a2_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001011000000100100000000000000100001000100011",
--  (1659) square_with_reduction_special_prime_2_16
-- reg_a = o1_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
"000110000001011000000000100000000000000100001000110111",
--  (1660) square_with_reduction_special_prime_2_17
-- -- In case of size 4
-- reg_a = a0_X; reg_b = a3_X; reg_acc = reg_o; o3_X = reg_o; Enable sign b; operation : 2*a*b + acc;
"000000100001011000010100100000000001010001101100000011",
--  (1661) square_with_reduction_special_prime_2_18
-- reg_a = a1_X; reg_b = a3_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001011000000100100000100001000100001100100011",
--  (1662) square_with_reduction_special_prime_2_19
-- reg_a = o1_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001011000000000100000000000000100001100110111",
--  (1663) square_with_reduction_special_prime_2_20
-- reg_a = a2_X; reg_b = a2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001011000000000100000000000000100001001000011",
--  (1664) square_with_reduction_special_prime_2_21
-- reg_a = o2_X; reg_b = primeSP2; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
"000000100001011000010000100000000000000100001001010111",
--  (1665) square_with_reduction_special_prime_2_22
-- reg_a = a2_X; reg_b = a3_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001011000000100100000100001000100001101000011",
--  (1666) square_with_reduction_special_prime_2_23
-- reg_a = o2_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001011000000000100000000000000100001101010111",
--  (1667) square_with_reduction_special_prime_2_24
-- reg_a = o3_X; reg_b = primeSP2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
"000000100001011000010000100000000000001000101001110111",
--  (1668) square_with_reduction_special_prime_2_25
-- reg_a = a3_X; reg_b = a3_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001011000000000100000100001100100001101100011",
--  (1669) square_with_reduction_special_prime_2_26
-- reg_a = o3_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; o3_X = reg_o >> 256; operation : a*b + acc;
"000000100001011001110000100000000000001101001101110111",
--  (1670) square_with_reduction_special_prime_2_27
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (1671) square_with_reduction_special_prime_2_28
-- -- In case of size 5, 6, 7, 8
-- reg_a = a0_X; reg_b = a3_X; reg_acc = reg_o; o3_X = reg_o; operation : 2*a*b + acc;
"000000100001100000010100100000000000010001101100000011",
--  (1672) square_with_reduction_special_prime_2_29
-- reg_a = o0_X; reg_b = primeSP4; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001100000000000100000100000000100010000010111",
--  (1673) square_with_reduction_special_prime_2_30
-- reg_a = a1_X; reg_b = a3_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001100000000100100000000000000100001100100011",
--  (1674) square_with_reduction_special_prime_2_31
-- reg_a = o1_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001100110111",
--  (1675) square_with_reduction_special_prime_2_32
-- reg_a = a2_X; reg_b = a2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001001000011",
--  (1676) square_with_reduction_special_prime_2_33
-- reg_a = o2_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
"001001000001100000000000100000000000000100001001010111",
--  (1677) square_with_reduction_special_prime_2_34
-- -- In case of size 5
-- reg_a = a0_X; reg_b = a4_X; reg_acc = reg_o; o4_X = reg_o; Enable sign b; operation : 2*a*b + acc;
"000000100001100000010100100000000001010110010000000011",
--  (1678) square_with_reduction_special_prime_2_35
-- reg_a = a1_X; reg_b = a4_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001100000000100100000100001000100010000100011",
--  (1679) square_with_reduction_special_prime_2_36
-- reg_a = o1_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100010000110111",
--  (1680) square_with_reduction_special_prime_2_37
-- reg_a = a2_X; reg_b = a3_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001100000000100100000000000000100001101000011",
--  (1681) square_with_reduction_special_prime_2_38
-- reg_a = o2_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001101010111",
--  (1682) square_with_reduction_special_prime_2_39
-- reg_a = o3_X; reg_b = primeSP2; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
"000000100001100000010000100000000000000100001001110111",
--  (1683) square_with_reduction_special_prime_2_40
-- reg_a = a2_X; reg_b = a4_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001100000000100100000100001000100010001000011",
--  (1684) square_with_reduction_special_prime_2_41
-- reg_a = o2_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100010001010111",
--  (1685) square_with_reduction_special_prime_2_42
-- reg_a = a3_X; reg_b = a3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001101100011",
--  (1686) square_with_reduction_special_prime_2_43
-- reg_a = o3_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001101110111",
--  (1687) square_with_reduction_special_prime_2_44
-- reg_a = o4_X; reg_b = primeSP2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
"000000100001100000010000100000000000001000101010010111",
--  (1688) square_with_reduction_special_prime_2_45
-- reg_a = a3_X; reg_b = a4_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001100000000100100000100001000100010001100011",
--  (1689) square_with_reduction_special_prime_2_46
-- reg_a = o3_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100010001110111",
--  (1690) square_with_reduction_special_prime_2_47
-- reg_a = o4_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
"000000100001100000010000100000000000001101001110010111",
--  (1691) square_with_reduction_special_prime_2_48
-- reg_a = a4_X; reg_b = a4_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001100000000000100000100001100100010010000011",
--  (1692) square_with_reduction_special_prime_2_49
-- reg_a = o4_X; reg_b = primeSP4; reg_acc = reg_o; o3_X = reg_o; o4_X = reg_o >> 256; operation : a*b + acc;
"000000100001100001110000100000000000010001110010010111",
--  (1693) square_with_reduction_special_prime_2_50
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (1694) square_with_reduction_special_prime_2_51
-- -- In case of sizes 6, 7, 8
-- reg_a = a0_X; reg_b = a4_X; reg_acc = reg_o; o4_X = reg_o; operation : 2*a*b + acc;
"000000100001101000010100100000000000010110010000000011",
--  (1695) square_with_reduction_special_prime_2_52
-- reg_a = o0_X; reg_b = primeSP5; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001101000000000100000100000000100010100010111",
--  (1696) square_with_reduction_special_prime_2_53
-- reg_a = a1_X; reg_b = a4_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001101000000100100000000000000100010000100011",
--  (1697) square_with_reduction_special_prime_2_54
-- reg_a = o1_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010000110111",
--  (1698) square_with_reduction_special_prime_2_55
-- reg_a = a2_X; reg_b = a3_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001101000000100100000000000000100001101000011",
--  (1699) square_with_reduction_special_prime_2_56
-- reg_a = o2_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001101010111",
--  (1700) square_with_reduction_special_prime_2_57
-- reg_a = o3_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
"001101000001101000000000100000000000000100001001110111",
--  (1701) square_with_reduction_special_prime_2_58
-- -- In case of size 6
-- reg_a = a0_X; reg_b = a5_X; reg_acc = reg_o; o5_X = reg_o; Enable sign b; operation : 2*a*b + acc;
"000000100001101000010100100000000001011010110100000011",
--  (1702) square_with_reduction_special_prime_2_59
-- reg_a = a1_X; reg_b = a5_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001101000000100100000100001000100010100100011",
--  (1703) square_with_reduction_special_prime_2_60
-- reg_a = o1_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010100110111",
--  (1704) square_with_reduction_special_prime_2_61
-- reg_a = a2_X; reg_b = a4_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001101000000100100000000000000100010001000011",
--  (1705) square_with_reduction_special_prime_2_62
-- reg_a = o2_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010001010111",
--  (1706) square_with_reduction_special_prime_2_63
-- reg_a = a3_X; reg_b = a3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001101100011",
--  (1707) square_with_reduction_special_prime_2_64
-- reg_a = o3_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001101110111",
--  (1708) square_with_reduction_special_prime_2_65
-- reg_a = o4_X; reg_b = primeSP2; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
"000000100001101000010000100000000000000100001010010111",
--  (1709) square_with_reduction_special_prime_2_66
-- reg_a = a2_X; reg_b = a5_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001101000000100100000100001000100010101000011",
--  (1710) square_with_reduction_special_prime_2_67
-- reg_a = o2_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010101010111",
--  (1711) square_with_reduction_special_prime_2_68
-- reg_a = a3_X; reg_b = a4_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001101000000100100000000000000100010001100011",
--  (1712) square_with_reduction_special_prime_2_69
-- reg_a = o3_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010001110111",
--  (1713) square_with_reduction_special_prime_2_70
-- reg_a = o4_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001110010111",
--  (1714) square_with_reduction_special_prime_2_71
-- reg_a = o5_X; reg_b = primeSP2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
"000000100001101000010000100000000000001000101010110111",
--  (1715) square_with_reduction_special_prime_2_72
-- reg_a = a3_X; reg_b = a5_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001101000000100100000100001000100010101100011",
--  (1716) square_with_reduction_special_prime_2_73
-- reg_a = o3_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010101110111",
--  (1717) square_with_reduction_special_prime_2_74
-- reg_a = a4_X; reg_b = a4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010010000011",
--  (1718) square_with_reduction_special_prime_2_75
-- reg_a = o4_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010010010111",
--  (1719) square_with_reduction_special_prime_2_76
-- reg_a = o5_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
"000000100001101000010000100000000000001101001110110111",
--  (1720) square_with_reduction_special_prime_2_77
-- reg_a = a4_X; reg_b = a5_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001101000000100100000100001000100010110000011",
--  (1721) square_with_reduction_special_prime_2_78
-- reg_a = o4_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010110010111",
--  (1722) square_with_reduction_special_prime_2_79
-- reg_a = o5_X; reg_b = primeSP4; reg_acc = reg_o; o3_X = reg_o; operation : a*b + acc;
"000000100001101000010000100000000000010001110010110111",
--  (1723) square_with_reduction_special_prime_2_80
-- reg_a = a5_X; reg_b = a5_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001101000000000100000100001100100010110100011",
--  (1724) square_with_reduction_special_prime_2_81
-- reg_a = o5_X; reg_b = primeSP5; reg_acc = reg_o; o4_X = reg_o; o5_X = reg_o >> 256; operation : a*b + acc;
"000000100001101001110000100000000000010110010110110111",
--  (1725) square_with_reduction_special_prime_2_82
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (1726) square_with_reduction_special_prime_2_83
-- -- In case of sizes 7, 8
-- reg_a = a0_X; reg_b = a5_X; reg_acc = reg_o; o5_X = reg_o; operation : 2*a*b + acc;
"000000100001110000010100100000000000011010110100000011",
--  (1727) square_with_reduction_special_prime_2_84
-- reg_a = o0_X; reg_b = primeSP6; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001110000000000100000100000000100011000010111",
--  (1728) square_with_reduction_special_prime_2_85
-- reg_a = a1_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001110000000100100000000000000100010100100011",
--  (1729) square_with_reduction_special_prime_2_86
-- reg_a = o1_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010100110111",
--  (1730) square_with_reduction_special_prime_2_87
-- reg_a = a2_X; reg_b = a4_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001110000000100100000000000000100010001000011",
--  (1731) square_with_reduction_special_prime_2_88
-- reg_a = o2_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010001010111",
--  (1732) square_with_reduction_special_prime_2_89
-- reg_a = a3_X; reg_b = a3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001101100011",
--  (1733) square_with_reduction_special_prime_2_90
-- reg_a = o3_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001101110111",
--  (1734) square_with_reduction_special_prime_2_91
-- reg_a = o4_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
"010001100001110000000000100000000000000100001010010111",
--  (1735) square_with_reduction_special_prime_2_92
-- -- In case of size 7
-- reg_a = a0_X; reg_b = a6_X; reg_acc = reg_o; o6_X = reg_o; Enable sign b; operation : 2*a*b + acc;
"000000100001110000010100100000000001011111011000000011",
--  (1736) square_with_reduction_special_prime_2_93
-- reg_a = a1_X; reg_b = a6_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001110000000100100000100001000100011000100011",
--  (1737) square_with_reduction_special_prime_2_94
-- reg_a = o1_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100011000110111",
--  (1738) square_with_reduction_special_prime_2_95
-- reg_a = a2_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001110000000100100000000000000100010101000011",
--  (1739) square_with_reduction_special_prime_2_96
-- reg_a = o2_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010101010111",
--  (1740) square_with_reduction_special_prime_2_97
-- reg_a = a3_X; reg_b = a4_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001110000000100100000000000000100010001100011",
--  (1741) square_with_reduction_special_prime_2_98
-- reg_a = o3_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010001110111",
--  (1742) square_with_reduction_special_prime_2_99
-- reg_a = o4_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001110010111",
--  (1743) square_with_reduction_special_prime_2_100
-- reg_a = o5_X; reg_b = primeSP2; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
"000000100001110000010000100000000000000100001010110111",
--  (1744) square_with_reduction_special_prime_2_101
-- reg_a = a2_X; reg_b = a6_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001110000000100100000100001000100011001000011",
--  (1745) square_with_reduction_special_prime_2_102
-- reg_a = o2_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100011001010111",
--  (1746) square_with_reduction_special_prime_2_103
-- reg_a = a3_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001110000000100100000000000000100010101100011",
--  (1747) square_with_reduction_special_prime_2_104
-- reg_a = o3_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010101110111",
--  (1748) square_with_reduction_special_prime_2_105
-- reg_a = a4_X; reg_b = a4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010010000011",
--  (1749) square_with_reduction_special_prime_2_106
-- reg_a = o4_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010010010111",
--  (1750) square_with_reduction_special_prime_2_107
-- reg_a = o5_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001110110111",
--  (1751) square_with_reduction_special_prime_2_108
-- reg_a = o6_X; reg_b = primeSP2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
"000000100001110000010000100000000000001000101011010111",
--  (1752) square_with_reduction_special_prime_2_109
-- reg_a = a3_X; reg_b = a6_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001110000000100100000100001000100011001100011",
--  (1753) square_with_reduction_special_prime_2_110
-- reg_a = o3_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100011001110111",
--  (1754) square_with_reduction_special_prime_2_111
-- reg_a = a4_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001110000000100100000000000000100010110000011",
--  (1755) square_with_reduction_special_prime_2_112
-- reg_a = o4_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010110010111",
--  (1756) square_with_reduction_special_prime_2_113
-- reg_a = o5_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010010110111",
--  (1757) square_with_reduction_special_prime_2_114
-- reg_a = o6_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
"000000100001110000010000100000000000001101001111010111",
--  (1758) square_with_reduction_special_prime_2_115
-- reg_a = a4_X; reg_b = a6_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001110000000100100000100001000100011010000011",
--  (1759) square_with_reduction_special_prime_2_116
-- reg_a = o4_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100011010010111",
--  (1760) square_with_reduction_special_prime_2_117
-- reg_a = a5_X; reg_b = a5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010110100011",
--  (1761) square_with_reduction_special_prime_2_118
-- reg_a = o5_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010110110111",
--  (1762) square_with_reduction_special_prime_2_119
-- reg_a = o6_X; reg_b = primeSP4; reg_acc = reg_o; o3_X = reg_o; operation : a*b + acc;
"000000100001110000010000100000000000010001110011010111",
--  (1763) square_with_reduction_special_prime_2_120
-- reg_a = a5_X; reg_b = a6_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001110000000100100000100001000100011010100011",
--  (1764) square_with_reduction_special_prime_2_121
-- reg_a = o5_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100011010110111",
--  (1765) square_with_reduction_special_prime_2_122
-- reg_a = o6_X; reg_b = primeSP5; reg_acc = reg_o; o4_X = reg_o; operation : a*b + acc;
"000000100001110000010000100000000000010110010111010111",
--  (1766) square_with_reduction_special_prime_2_123
-- reg_a = a6_X; reg_b = a6_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001110000000000100000100001100100011011000011",
--  (1767) square_with_reduction_special_prime_2_124
-- reg_a = o6_X; reg_b = primeSP6; reg_acc = reg_o; o5_X = reg_o; o6_X = reg_o >> 256; operation : a*b + acc;
"000000100001110001110000100000000000011010111011010111",
--  (1768) square_with_reduction_special_prime_2_125
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (1769) square_with_reduction_special_prime_2_126
-- -- In case of size 8
-- reg_a = a0_X; reg_b = a6_X; reg_acc = reg_o; o6_X = reg_o; operation : 2*a*b + acc;
"000000100001111000010100100000000000011111011000000011",
--  (1770) square_with_reduction_special_prime_2_127
-- reg_a = o0_X; reg_b = primeSP7; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001111000000000100000100000000100011100010111",
--  (1771) square_with_reduction_special_prime_2_128
-- reg_a = a1_X; reg_b = a6_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001111000000100100000000000000100011000100011",
--  (1772) square_with_reduction_special_prime_2_129
-- reg_a = o1_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011000110111",
--  (1773) square_with_reduction_special_prime_2_130
-- reg_a = a2_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001111000000100100000000000000100010101000011",
--  (1774) square_with_reduction_special_prime_2_131
-- reg_a = o2_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010101010111",
--  (1775) square_with_reduction_special_prime_2_132
-- reg_a = a3_X; reg_b = a4_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001111000000100100000000000000100010001100011",
--  (1776) square_with_reduction_special_prime_2_133
-- reg_a = o3_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010001110111",
--  (1777) square_with_reduction_special_prime_2_134
-- reg_a = o4_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001110010111",
--  (1778) square_with_reduction_special_prime_2_135
-- reg_a = o5_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001010110111",
--  (1779) square_with_reduction_special_prime_2_136
-- reg_a = a0_X; reg_b = a7_X; reg_acc = reg_o; o7_X = reg_o; Enable sign b; operation : 2*a*b + acc;
"000000100001111000010100100000000001000011111100000011",
--  (1780) square_with_reduction_special_prime_2_137
-- reg_a = a1_X; reg_b = a7_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001111000000100100000100001000100011100100011",
--  (1781) square_with_reduction_special_prime_2_138
-- reg_a = o1_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011100110111",
--  (1782) square_with_reduction_special_prime_2_139
-- reg_a = a2_X; reg_b = a6_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001111000000100100000000000000100011001000011",
--  (1783) square_with_reduction_special_prime_2_140
-- reg_a = o2_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011001010111",
--  (1784) square_with_reduction_special_prime_2_141
-- reg_a = a3_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001111000000100100000000000000100010101100011",
--  (1785) square_with_reduction_special_prime_2_142
-- reg_a = o3_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010101110111",
--  (1786) square_with_reduction_special_prime_2_143
-- reg_a = a4_X; reg_b = a4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010010000011",
--  (1787) square_with_reduction_special_prime_2_144
-- reg_a = o4_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010010010111",
--  (1788) square_with_reduction_special_prime_2_145
-- reg_a = o5_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001110110111",
--  (1789) square_with_reduction_special_prime_2_146
-- reg_a = o6_X; reg_b = primeSP2; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000000100001011010111",
--  (1790) square_with_reduction_special_prime_2_147
-- reg_a = a2_X; reg_b = a7_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001111000000100100000100001000100011101000011",
--  (1791) square_with_reduction_special_prime_2_148
-- reg_a = o2_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011101010111",
--  (1792) square_with_reduction_special_prime_2_149
-- reg_a = a3_X; reg_b = a6_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001111000000100100000000000000100011001100011",
--  (1793) square_with_reduction_special_prime_2_150
-- reg_a = o3_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011001110111",
--  (1794) square_with_reduction_special_prime_2_151
-- reg_a = a4_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001111000000100100000000000000100010110000011",
--  (1795) square_with_reduction_special_prime_2_152
-- reg_a = o4_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010110010111",
--  (1796) square_with_reduction_special_prime_2_153
-- reg_a = o5_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010010110111",
--  (1797) square_with_reduction_special_prime_2_154
-- reg_a = o6_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001111010111",
--  (1798) square_with_reduction_special_prime_2_155
-- reg_a = o7_X; reg_b = primeSP2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000001000101011110111",
--  (1799) square_with_reduction_special_prime_2_156
-- reg_a = a3_X; reg_b = a7_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001111000000100100000100001000100011101100011",
--  (1800) square_with_reduction_special_prime_2_157
-- reg_a = o3_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011101110111",
--  (1801) square_with_reduction_special_prime_2_158
-- reg_a = a4_X; reg_b = a6_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001111000000100100000000000000100011010000011",
--  (1802) square_with_reduction_special_prime_2_159
-- reg_a = o4_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011010010111",
--  (1803) square_with_reduction_special_prime_2_160
-- reg_a = a5_X; reg_b = a5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010110100011",
--  (1804) square_with_reduction_special_prime_2_161
-- reg_a = o5_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010110110111",
--  (1805) square_with_reduction_special_prime_2_162
-- reg_a = o6_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010011010111",
--  (1806) square_with_reduction_special_prime_2_163
-- reg_a = o7_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000001101001111110111",
--  (1807) square_with_reduction_special_prime_2_164
-- reg_a = a4_X; reg_b = a7_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001111000000100100000100001000100011110000011",
--  (1808) square_with_reduction_special_prime_2_165
-- reg_a = o4_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011110010111",
--  (1809) square_with_reduction_special_prime_2_166
-- reg_a = a5_X; reg_b = a6_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001111000000100100000000000000100011010100011",
--  (1810) square_with_reduction_special_prime_2_167
-- reg_a = o5_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011010110111",
--  (1811) square_with_reduction_special_prime_2_168
-- reg_a = o6_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010111010111",
--  (1812) square_with_reduction_special_prime_2_169
-- reg_a = o7_X; reg_b = primeSP4; reg_acc = reg_o; o3_X = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000010001110011110111",
--  (1813) square_with_reduction_special_prime_2_170
-- reg_a = a5_X; reg_b = a7_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001111000000100100000100001000100011110100011",
--  (1814) square_with_reduction_special_prime_2_171
-- reg_a = o5_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011110110111",
--  (1815) square_with_reduction_special_prime_2_172
-- reg_a = a6_X; reg_b = a6_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011011000011",
--  (1816) square_with_reduction_special_prime_2_173
-- reg_a = o6_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011011010111",
--  (1817) square_with_reduction_special_prime_2_174
-- reg_a = o7_X; reg_b = primeSP5; reg_acc = reg_o; o4_X = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000010110010111110111",
--  (1818) square_with_reduction_special_prime_2_175
-- reg_a = a6_X; reg_b = a7_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001111000000100100000100001000100011111000011",
--  (1819) square_with_reduction_special_prime_2_176
-- reg_a = o6_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011111010111",
--  (1820) square_with_reduction_special_prime_2_177
-- reg_a = o7_X; reg_b = primeSP6; reg_acc = reg_o; o5_X = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000011010111011110111",
--  (1821) square_with_reduction_special_prime_2_178
-- reg_a = a7_X; reg_b = a7_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001111000000000100000100001100100011111100011",
--  (1822) square_with_reduction_special_prime_2_179
-- reg_a = o7_X; reg_b = primeSP7; reg_acc = reg_o; o6_X = reg_o; o7_X = reg_o >> 256; operation : a*b + acc;
"000000100001111001110000100000000000011111011111110111",
--  (1823) square_with_reduction_special_prime_2_180
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (1824) square_with_reduction_special_prime_3_0
-- -- In case of sizes 3, 4, 5, 6, 7, 8
-- reg_a = a0_X; reg_b = a0_X; reg_acc = 0; o0_X = reg_o; operation : a*b + acc;
"000000100001010000010000100000010000000100000000000011",
--  (1825) square_with_reduction_special_prime_3_1
-- reg_a = a0_X; reg_b = a1_X; reg_acc = reg_o >> 256; o1_X = reg_o; operation : 2*a*b + acc;
"000000100001010000010100100000100000001000100100000011",
--  (1826) square_with_reduction_special_prime_3_2
-- reg_a = a1_X; reg_b = a1_X; reg_acc = reg_o >> 256; operation : a*b + acc;
"000010100001010000000000100000100000000100000100100011",
--  (1827) square_with_reduction_special_prime_3_3
-- -- In case of size 3
-- reg_a = a0_X; reg_b = a2_X; reg_acc = reg_o; o2_X = reg_o; Enable sign b; operation : 2*a*b + acc;
"000000100001010000010100100000000001001101001000000011",
--  (1828) square_with_reduction_special_prime_3_4
-- reg_a = a1_X; reg_b = a2_X; reg_acc = reg_o >> 256; Enable sign b; o0_X = reg_o; operation : 2*a*b + acc;
"000000100001010000010100100000100001000100001000100011",
--  (1829) square_with_reduction_special_prime_3_5
-- reg_a = a2_X; reg_b = a2_X; reg_acc = reg_o >> 256; Enable sign a,b; o1_X = reg_o; o2_X = reg_o >> 256; operation : a*b + acc;
"000000100001010001110000100000100001101000101001000011",
--  (1830) square_with_reduction_special_prime_3_6
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (1831) square_with_reduction_special_prime_3_7
-- -- In case of sizes 4, 5, 6, 7, 8
-- reg_a = a0_X; reg_b = a2_X; reg_acc = reg_o; o2_X = reg_o; operation : 2*a*b + acc;
"000000100001011000010100100000000000001101001000000011",
--  (1832) square_with_reduction_special_prime_3_8
-- reg_a = o0_X; reg_b = primeSP3; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001011000000000100000100000000100001100010111",
--  (1833) square_with_reduction_special_prime_3_9
-- reg_a = a1_X; reg_b = a2_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000101000001011000000100100000000000000100001000100011",
--  (1834) square_with_reduction_special_prime_3_10
-- -- In case of size 4
-- reg_a = a0_X; reg_b = a3_X; reg_acc = reg_o; o3_X = reg_o; Enable sign b; operation : 2*a*b + acc;
"000000100001011000010100100000000001010001101100000011",
--  (1835) square_with_reduction_special_prime_3_11
-- reg_a = a1_X; reg_b = a3_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001011000000100100000100001000100001100100011",
--  (1836) square_with_reduction_special_prime_3_12
-- reg_a = o1_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001011000000000100000000000000100001100110111",
--  (1837) square_with_reduction_special_prime_3_13
-- reg_a = a2_X; reg_b = a2_X; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
"000000100001011000010000100000000000000100001001000011",
--  (1838) square_with_reduction_special_prime_3_14
-- reg_a = a2_X; reg_b = a3_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001011000000100100000100001000100001101000011",
--  (1839) square_with_reduction_special_prime_3_15
-- reg_a = o2_X; reg_b = primeSP3; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
"000000100001011000010000100000000000001000101101010111",
--  (1840) square_with_reduction_special_prime_3_16
-- reg_a = a3_X; reg_b = a3_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001011000000000100000100001100100001101100011",
--  (1841) square_with_reduction_special_prime_3_17
-- reg_a = o3_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; o3_X = reg_o >> 256; operation : a*b + acc;
"000000100001011001110000100000000000001101001101110111",
--  (1842) square_with_reduction_special_prime_3_18
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (1843) square_with_reduction_special_prime_3_19
-- -- In case of sizes 5, 6, 7, 8
-- reg_a = a0_X; reg_b = a3_X; reg_acc = reg_o; o3_X = reg_o; operation : 2*a*b + acc;
"000000100001100000010100100000000000010001101100000011",
--  (1844) square_with_reduction_special_prime_3_20
-- reg_a = o0_X; reg_b = primeSP4; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001100000000000100000100000000100010000010111",
--  (1845) square_with_reduction_special_prime_3_21
-- reg_a = a1_X; reg_b = a3_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001100000000100100000000000000100001100100011",
--  (1846) square_with_reduction_special_prime_3_22
-- reg_a = o1_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001100110111",
--  (1847) square_with_reduction_special_prime_3_23
-- reg_a = a2_X; reg_b = a2_X; reg_acc = reg_o; operation : a*b + acc;
"001000000001100000000000100000000000000100001001000011",
--  (1848) square_with_reduction_special_prime_3_24
-- -- In case of size 5
-- reg_a = a0_X; reg_b = a4_X; reg_acc = reg_o; o4_X = reg_o; Enable sign b; operation : 2*a*b + acc;
"000000100001100000010100100000000001010110010000000011",
--  (1849) square_with_reduction_special_prime_3_25
-- reg_a = a1_X; reg_b = a4_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001100000000100100000100001000100010000100011",
--  (1850) square_with_reduction_special_prime_3_26
-- reg_a = o1_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100010000110111",
--  (1851) square_with_reduction_special_prime_3_27
-- reg_a = a2_X; reg_b = a3_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001100000000100100000000000000100001101000011",
--  (1852) square_with_reduction_special_prime_3_28
-- reg_a = o2_X; reg_b = primeSP3; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
"000000100001100000010000100000000000000100001101010111",
--  (1853) square_with_reduction_special_prime_3_29
-- reg_a = a2_X; reg_b = a4_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001100000000100100000100001000100010001000011",
--  (1854) square_with_reduction_special_prime_3_30
-- reg_a = o2_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100010001010111",
--  (1855) square_with_reduction_special_prime_3_31
-- reg_a = a3_X; reg_b = a3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001101100011",
--  (1856) square_with_reduction_special_prime_3_32
-- reg_a = o3_X; reg_b = primeSP3; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
"000000100001100000010000100000000000001000101101110111",
--  (1857) square_with_reduction_special_prime_3_33
-- reg_a = a3_X; reg_b = a4_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001100000000100100000100001000100010001100011",
--  (1858) square_with_reduction_special_prime_3_34
-- reg_a = o3_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100010001110111",
--  (1859) square_with_reduction_special_prime_3_35
-- reg_a = o4_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
"000000100001100000010000100000000000001101001110010111",
--  (1860) square_with_reduction_special_prime_3_36
-- reg_a = a4_X; reg_b = a4_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001100000000000100000100001100100010010000011",
--  (1861) square_with_reduction_special_prime_3_37
-- reg_a = o4_X; reg_b = primeSP4; reg_acc = reg_o; o3_X = reg_o; o4_X = reg_o >> 256; operation : a*b + acc;
"000000100001100001110000100000000000010001110010010111",
--  (1862) square_with_reduction_special_prime_3_38
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (1863) square_with_reduction_special_prime_3_39
-- -- In case of sizes 6, 7, 8
-- reg_a = a0_X; reg_b = a4_X; reg_acc = reg_o; o4_X = reg_o; operation : 2*a*b + acc;
"000000100001101000010100100000000000010110010000000011",
--  (1864) square_with_reduction_special_prime_3_40
-- reg_a = o0_X; reg_b = primeSP5; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001101000000000100000100000000100010100010111",
--  (1865) square_with_reduction_special_prime_3_41
-- reg_a = a1_X; reg_b = a4_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001101000000100100000000000000100010000100011",
--  (1866) square_with_reduction_special_prime_3_42
-- reg_a = o1_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010000110111",
--  (1867) square_with_reduction_special_prime_3_43
-- reg_a = a2_X; reg_b = a3_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001101000000100100000000000000100001101000011",
--  (1868) square_with_reduction_special_prime_3_44
-- reg_a = o2_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"001100000001101000000000100000000000000100001101010111",
--  (1869) square_with_reduction_special_prime_3_45
-- -- In case of size 6
-- reg_a = a0_X; reg_b = a5_X; reg_acc = reg_o; o5_X = reg_o; Enable sign b; operation : 2*a*b + acc;
"000000100001101000010100100000000001011010110100000011",
--  (1870) square_with_reduction_special_prime_3_46
-- reg_a = a1_X; reg_b = a5_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001101000000100100000100001000100010100100011",
--  (1871) square_with_reduction_special_prime_3_47
-- reg_a = o1_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010100110111",
--  (1872) square_with_reduction_special_prime_3_48
-- reg_a = a2_X; reg_b = a4_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001101000000100100000000000000100010001000011",
--  (1873) square_with_reduction_special_prime_3_49
-- reg_a = o2_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010001010111",
--  (1874) square_with_reduction_special_prime_3_50
-- reg_a = a3_X; reg_b = a3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001101100011",
--  (1875) square_with_reduction_special_prime_3_51
-- reg_a = o3_X; reg_b = primeSP3; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
"000000100001101000010000100000000000000100001101110111",
--  (1876) square_with_reduction_special_prime_3_52
-- reg_a = a2_X; reg_b = a5_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001101000000100100000100001000100010101000011",
--  (1877) square_with_reduction_special_prime_3_53
-- reg_a = o2_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010101010111",
--  (1878) square_with_reduction_special_prime_3_54
-- reg_a = a3_X; reg_b = a4_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001101000000100100000000000000100010001100011",
--  (1879) square_with_reduction_special_prime_3_55
-- reg_a = o3_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010001110111",
--  (1880) square_with_reduction_special_prime_3_56
-- reg_a = o4_X; reg_b = primeSP3; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
"000000100001101000010000100000000000001000101110010111",
--  (1881) square_with_reduction_special_prime_3_57
-- reg_a = a3_X; reg_b = a5_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001101000000100100000100001000100010101100011",
--  (1882) square_with_reduction_special_prime_3_58
-- reg_a = o3_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010101110111",
--  (1883) square_with_reduction_special_prime_3_59
-- reg_a = a4_X; reg_b = a4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010010000011",
--  (1884) square_with_reduction_special_prime_3_60
-- reg_a = o4_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010010010111",
--  (1885) square_with_reduction_special_prime_3_61
-- reg_a = o5_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
"000000100001101000010000100000000000001101001110110111",
--  (1886) square_with_reduction_special_prime_3_62
-- reg_a = a4_X; reg_b = a5_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001101000000100100000100001000100010110000011",
--  (1887) square_with_reduction_special_prime_3_63
-- reg_a = o4_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010110010111",
--  (1888) square_with_reduction_special_prime_3_64
-- reg_a = o5_X; reg_b = primeSP4; reg_acc = reg_o; o3_X = reg_o; operation : a*b + acc;
"000000100001101000010000100000000000010001110010110111",
--  (1889) square_with_reduction_special_prime_3_65
-- reg_a = a5_X; reg_b = a5_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001101000000000100000100001100100010110100011",
--  (1890) square_with_reduction_special_prime_3_66
-- reg_a = o5_X; reg_b = primeSP5; reg_acc = reg_o; o4_X = reg_o; o5_X = reg_o >> 256; operation : a*b + acc;
"000000100001101001110000100000000000010110010110110111",
--  (1891) square_with_reduction_special_prime_3_67
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (1892) square_with_reduction_special_prime_3_68
-- -- In case of sizes 7, 8
-- reg_a = a0_X; reg_b = a5_X; reg_acc = reg_o; o5_X = reg_o; operation : 2*a*b + acc;
"000000100001110000010100100000000000011010110100000011",
--  (1893) square_with_reduction_special_prime_3_69
-- reg_a = o0_X; reg_b = primeSP6; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001110000000000100000100000000100011000010111",
--  (1894) square_with_reduction_special_prime_3_70
-- reg_a = a1_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001110000000100100000000000000100010100100011",
--  (1895) square_with_reduction_special_prime_3_71
-- reg_a = o1_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010100110111",
--  (1896) square_with_reduction_special_prime_3_72
-- reg_a = a2_X; reg_b = a4_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001110000000100100000000000000100010001000011",
--  (1897) square_with_reduction_special_prime_3_73
-- reg_a = o2_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010001010111",
--  (1898) square_with_reduction_special_prime_3_74
-- reg_a = a3_X; reg_b = a3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001101100011",
--  (1899) square_with_reduction_special_prime_3_75
-- reg_a = o3_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"010000100001110000000000100000000000000100001101110111",
--  (1900) square_with_reduction_special_prime_3_76
-- -- In case of size 7
-- reg_a = a0_X; reg_b = a6_X; reg_acc = reg_o; o6_X = reg_o; Enable sign b; operation : 2*a*b + acc;
"000000100001110000010100100000000001011111011000000011",
--  (1901) square_with_reduction_special_prime_3_77
-- reg_a = a1_X; reg_b = a6_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001110000000100100000100001000100011000100011",
--  (1902) square_with_reduction_special_prime_3_78
-- reg_a = o1_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100011000110111",
--  (1903) square_with_reduction_special_prime_3_79
-- reg_a = a2_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001110000000100100000000000000100010101000011",
--  (1904) square_with_reduction_special_prime_3_80
-- reg_a = o2_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010101010111",
--  (1905) square_with_reduction_special_prime_3_81
-- reg_a = a3_X; reg_b = a4_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001110000000100100000000000000100010001100011",
--  (1906) square_with_reduction_special_prime_3_82
-- reg_a = o3_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010001110111",
--  (1907) square_with_reduction_special_prime_3_83
-- reg_a = o4_X; reg_b = primeSP3; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
"000000100001110000010000100000000000000100001110010111",
--  (1908) square_with_reduction_special_prime_3_84
-- reg_a = a2_X; reg_b = a6_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001110000000100100000100001000100011001000011",
--  (1909) square_with_reduction_special_prime_3_85
-- reg_a = o2_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100011001010111",
--  (1910) square_with_reduction_special_prime_3_86
-- reg_a = a3_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001110000000100100000000000000100010101100011",
--  (1911) square_with_reduction_special_prime_3_87
-- reg_a = o3_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010101110111",
--  (1912) square_with_reduction_special_prime_3_88
-- reg_a = a4_X; reg_b = a4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010010000011",
--  (1913) square_with_reduction_special_prime_3_89
-- reg_a = o4_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010010010111",
--  (1914) square_with_reduction_special_prime_3_90
-- reg_a = o5_X; reg_b = primeSP3; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
"000000100001110000010000100000000000001000101110110111",
--  (1915) square_with_reduction_special_prime_3_91
-- reg_a = a3_X; reg_b = a6_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001110000000100100000100001000100011001100011",
--  (1916) square_with_reduction_special_prime_3_92
-- reg_a = o3_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100011001110111",
--  (1917) square_with_reduction_special_prime_3_93
-- reg_a = a4_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001110000000100100000000000000100010110000011",
--  (1918) square_with_reduction_special_prime_3_94
-- reg_a = o4_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010110010111",
--  (1919) square_with_reduction_special_prime_3_95
-- reg_a = o5_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010010110111",
--  (1920) square_with_reduction_special_prime_3_96
-- reg_a = o6_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
"000000100001110000010000100000000000001101001111010111",
--  (1921) square_with_reduction_special_prime_3_97
-- reg_a = a4_X; reg_b = a6_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001110000000100100000100001000100011010000011",
--  (1922) square_with_reduction_special_prime_3_98
-- reg_a = o4_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100011010010111",
--  (1923) square_with_reduction_special_prime_3_99
-- reg_a = a5_X; reg_b = a5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010110100011",
--  (1924) square_with_reduction_special_prime_3_100
-- reg_a = o5_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010110110111",
--  (1925) square_with_reduction_special_prime_3_101
-- reg_a = o6_X; reg_b = primeSP4; reg_acc = reg_o; o3_X = reg_o; operation : a*b + acc;
"000000100001110000010000100000000000010001110011010111",
--  (1926) square_with_reduction_special_prime_3_102
-- reg_a = a5_X; reg_b = a6_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001110000000100100000100001000100011010100011",
--  (1927) square_with_reduction_special_prime_3_103
-- reg_a = o5_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100011010110111",
--  (1928) square_with_reduction_special_prime_3_104
-- reg_a = o6_X; reg_b = primeSP5; reg_acc = reg_o; o4_X = reg_o; operation : a*b + acc;
"000000100001110000010000100000000000010110010111010111",
--  (1929) square_with_reduction_special_prime_3_105
-- reg_a = a6_X; reg_b = a6_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001110000000000100000100001100100011011000011",
--  (1930) square_with_reduction_special_prime_3_106
-- reg_a = o6_X; reg_b = primeSP6; reg_acc = reg_o; o5_X = reg_o; o6_X = reg_o >> 256; operation : a*b + acc;
"000000100001110001110000100000000000011010111011010111",
--  (1931) square_with_reduction_special_prime_3_107
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (1932) square_with_reduction_special_prime_3_108
-- -- In case of size 8
-- reg_a = a0_X; reg_b = a6_X; reg_acc = reg_o; o6_X = reg_o; operation : 2*a*b + acc;
"000000100001111000010100100000000000011011011000000011",
--  (1933) square_with_reduction_special_prime_3_109
-- reg_a = o0_X; reg_b = primeSP7; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001111000000000100000100000000100011100010111",
--  (1934) square_with_reduction_special_prime_3_110
-- reg_a = a1_X; reg_b = a6_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001111000000100100000000000000100011000100011",
--  (1935) square_with_reduction_special_prime_3_111
-- reg_a = o1_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011000110111",
--  (1936) square_with_reduction_special_prime_3_112
-- reg_a = a2_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001111000000100100000000000000100010101000011",
--  (1937) square_with_reduction_special_prime_3_113
-- reg_a = o2_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010101010111",
--  (1938) square_with_reduction_special_prime_3_114
-- reg_a = a3_X; reg_b = a4_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001111000000100100000000000000100010001100011",
--  (1939) square_with_reduction_special_prime_3_115
-- reg_a = o3_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010001110111",
--  (1940) square_with_reduction_special_prime_3_116
-- reg_a = o4_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001110010111",
--  (1941) square_with_reduction_special_prime_3_117
-- reg_a = a0_X; reg_b = a7_X; reg_acc = reg_o; o7_X = reg_o; Enable sign b; operation : 2*a*b + acc;
"000000100001111000010100100000000001011111111100000011",
--  (1942) square_with_reduction_special_prime_3_118
-- reg_a = a1_X; reg_b = a7_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001111000000100100000100001000100011100100011",
--  (1943) square_with_reduction_special_prime_3_119
-- reg_a = o1_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011100110111",
--  (1944) square_with_reduction_special_prime_3_120
-- reg_a = a2_X; reg_b = a6_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001111000000100100000000000000100011001000011",
--  (1945) square_with_reduction_special_prime_3_121
-- reg_a = o2_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011001010111",
--  (1946) square_with_reduction_special_prime_3_122
-- reg_a = a3_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001111000000100100000000000000100010101100011",
--  (1947) square_with_reduction_special_prime_3_123
-- reg_a = o3_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010101110111",
--  (1948) square_with_reduction_special_prime_3_124
-- reg_a = a4_X; reg_b = a4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010010000011",
--  (1949) square_with_reduction_special_prime_3_125
-- reg_a = o4_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010010010111",
--  (1950) square_with_reduction_special_prime_3_126
-- reg_a = o5_X; reg_b = primeSP3; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000000100001110110111",
--  (1951) square_with_reduction_special_prime_3_127
-- reg_a = a2_X; reg_b = a7_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001111000000100100000100001000100011101000011",
--  (1952) square_with_reduction_special_prime_3_128
-- reg_a = o2_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011101010111",
--  (1953) square_with_reduction_special_prime_3_129
-- reg_a = a3_X; reg_b = a6_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001111000000100100000000000000100011001100011",
--  (1954) square_with_reduction_special_prime_3_130
-- reg_a = o3_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011001110111",
--  (1955) square_with_reduction_special_prime_3_131
-- reg_a = a4_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001111000000100100000000000000100010110000011",
--  (1956) square_with_reduction_special_prime_3_132
-- reg_a = o4_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010110010111",
--  (1957) square_with_reduction_special_prime_3_133
-- reg_a = o5_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010010110111",
--  (1958) square_with_reduction_special_prime_3_134
-- reg_a = o6_X; reg_b = primeSP3; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000001000101111010111",
--  (1959) square_with_reduction_special_prime_3_135
-- reg_a = a3_X; reg_b = a7_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001111000000100100000100001000100011101100011",
--  (1960) square_with_reduction_special_prime_3_136
-- reg_a = o3_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011101110111",
--  (1961) square_with_reduction_special_prime_3_137
-- reg_a = a4_X; reg_b = a6_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001111000000100100000000000000100011010000011",
--  (1962) square_with_reduction_special_prime_3_138
-- reg_a = o4_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011010010111",
--  (1963) square_with_reduction_special_prime_3_139
-- reg_a = a5_X; reg_b = a5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010110100011",
--  (1964) square_with_reduction_special_prime_3_140
-- reg_a = o5_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010110110111",
--  (1965) square_with_reduction_special_prime_3_141
-- reg_a = o6_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010011010111",
--  (1966) square_with_reduction_special_prime_3_142
-- reg_a = o7_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000001101001111110111",
--  (1967) square_with_reduction_special_prime_3_143
-- reg_a = a4_X; reg_b = a7_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001111000000100100000100001000100011110000011",
--  (1968) square_with_reduction_special_prime_3_144
-- reg_a = o4_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011110010111",
--  (1969) square_with_reduction_special_prime_3_145
-- reg_a = a5_X; reg_b = a6_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001111000000100100000000000000100011010100011",
--  (1970) square_with_reduction_special_prime_3_146
-- reg_a = o5_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011010110111",
--  (1971) square_with_reduction_special_prime_3_147
-- reg_a = o6_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010111010111",
--  (1972) square_with_reduction_special_prime_3_148
-- reg_a = o7_X; reg_b = primeSP4; reg_acc = reg_o; o3_X = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000010001110011110111",
--  (1973) square_with_reduction_special_prime_3_149
-- reg_a = a5_X; reg_b = a7_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001111000000100100000100001000100011110100011",
--  (1974) square_with_reduction_special_prime_3_150
-- reg_a = o5_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011110110111",
--  (1975) square_with_reduction_special_prime_3_151
-- reg_a = a6_X; reg_b = a6_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011011000011",
--  (1976) square_with_reduction_special_prime_3_152
-- reg_a = o6_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011011010111",
--  (1977) square_with_reduction_special_prime_3_153
-- reg_a = o7_X; reg_b = primeSP5; reg_acc = reg_o; o4_X = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000010110010111110111",
--  (1978) square_with_reduction_special_prime_3_154
-- reg_a = a6_X; reg_b = a7_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001111000000100100000100001000100011111000011",
--  (1979) square_with_reduction_special_prime_3_155
-- reg_a = o6_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011111010111",
--  (1980) square_with_reduction_special_prime_3_156
-- reg_a = o7_X; reg_b = primeSP6; reg_acc = reg_o; o5_X = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000011010111011110111",
--  (1981) square_with_reduction_special_prime_3_157
-- reg_a = a7_X; reg_b = a7_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001111000000000100000100001100100011111100011",
--  (1982) square_with_reduction_special_prime_3_158
-- reg_a = o7_X; reg_b = primeSP7; reg_acc = reg_o; o6_X = reg_o; o7_X = reg_o >> 256; operation : a*b + acc;
"000000100001111001110000100000000000011111011111110111",
--  (1983) square_with_reduction_special_prime_3_159
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (1984) addition_subtraction_direct_0
-- -- In case of size 1
-- reg_a = a0_X; reg_b = b0_X; reg_acc = 0; o0_0 = reg_o; Enable sign a,b; operation : b +/- a + acc;
"000000100001000000010000001000010001100100000000000010",
--  (1985) addition_subtraction_direct_1
-- NOP 4 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : b + a + acc;
"000000000000000100000000010000011110000100000000000010",
--  (1986) addition_subtraction_direct_2
-- -- In case of size 2, 3, 4, 5, 6, 7, 8
-- reg_a = a0_X; reg_b = b0_X; reg_acc = 0; o0_X = reg_o; operation : b +/- a + acc;
"000001100001001000010000001000010000000100000000000010",
--  (1987) addition_subtraction_direct_3
-- -- In case of size 2
-- reg_a = a1_X; reg_b = b1_X; reg_acc = reg_o >> 256; o1_X = reg_o; Enable sign a, b; operation : b +/- a + acc;
"000000100001001000010000001000100001101000100100100010",
--  (1988) addition_subtraction_direct_4
-- NOP 4 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : b + a + acc;
"000000000000000100000000010000011110000100000000000010",
--  (1989) addition_subtraction_direct_5
-- -- In case of size 3, 4, 5, 6, 7, 8
-- reg_a = a1_X; reg_b = b1_X; reg_acc = reg_o >> 256; o1_X = reg_o; operation : b +/- a + acc;
"000001100001010000010000001000100000001000100100100010",
--  (1990) addition_subtraction_direct_6
-- -- In case of size 3
-- reg_a = a2_X; reg_b = b2_X; reg_acc = reg_o >> 256; o2_X = reg_o; Enable sign a,b; operation : b +/- a + acc;
"000000100001010000010000001000100001100101001001000010",
--  (1991) addition_subtraction_direct_7
-- NOP 4 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : b + a + acc;
"000000000000000100000000010000011110000100000000000010",
--  (1992) addition_subtraction_direct_8
-- -- In case of size 4, 5, 6, 7, 8
-- reg_a = a2_X; reg_b = b2_X; reg_acc = reg_o >> 256; o2_X = reg_o; operation : b +/- a + acc;
"000001100001011000010000001000100000000101001001000010",
--  (1993) addition_subtraction_direct_9
-- -- In case of size 4
-- reg_a = a3_X; reg_b = b3_X; reg_acc = reg_o >> 256; o3_X = reg_o; Enable sign a,b; operation : b +/- a + acc;
"000000100001011000010000001000100001110001101101100010",
--  (1994) addition_subtraction_direct_10
-- NOP 4 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : b + a + acc;
"000000000000000100000000010000011110000100000000000010",
--  (1995) addition_subtraction_direct_11
-- -- In case of size 4, 5, 6, 7, 8
-- reg_a = a3_X; reg_b = b3_X; reg_acc = reg_o >> 256; o3_X = reg_o; operation : b +/- a + acc;
"000001100001100000010000001000100000010001101101100010",
--  (1996) addition_subtraction_direct_12
-- -- In case of size 5
-- reg_a = a4_X; reg_b = b4_X; reg_acc = reg_o >> 256; o4_X = reg_o; Enable sign a,b; operation : b +/- a + acc;
"000000100001100000010000001000100001110110010010000010",
--  (1997) addition_subtraction_direct_13
-- NOP 4 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : b + a + acc;
"000000000000000100000000010000011110000100000000000010",
--  (1998) addition_subtraction_direct_14
-- -- In case of size 6, 7, 8
-- reg_a = a4_X; reg_b = b4_X; reg_acc = reg_o >> 256; o4_X = reg_o; operation : b +/- a + acc;
"000001100001101000010000001000100000010110010010000010",
--  (1999) addition_subtraction_direct_15
-- -- In case of size 6
-- reg_a = a5_X; reg_b = b5_X; reg_acc = reg_o >> 256; o5_X = reg_o; Enable sign a,b; operation : b +/- a + acc;
"000000100001101000010000001000100001111010110110100010",
--  (2000) addition_subtraction_direct_16
-- NOP 4 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : b + a + acc;
"000000000000000100000000010000011110000100000000000010",
--  (2001) addition_subtraction_direct_17
-- -- In case of size 7, 8
-- reg_a = a5_X; reg_b = b5_X; reg_acc = reg_o >> 256; o5_X = reg_o; operation : b +/- a + acc;
"000001100001110000010000001000100000011010110110100010",
--  (2002) addition_subtraction_direct_18
-- -- In case of size 7
-- reg_a = a6_X; reg_b = b6_X; reg_acc = reg_o >> 256; o6_X = reg_o; Enable sign a,b; operation : b +/- a + acc;
"000000100001110000010000001000100001111111011011000010",
--  (2003) addition_subtraction_direct_19
-- NOP 4 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : b + a + acc;
"000000000000000100000000010000011110000100000000000010",
--  (2004) addition_subtraction_direct_20
-- -- In case of size 8
-- reg_a = a6_X; reg_b = b6_X; reg_acc = reg_o >> 256; o6_X = reg_o; operation : b +/- a + acc;
"000000100001111000010000001000100000011111011011000010",
--  (2005) addition_subtraction_direct_21
-- reg_a = a7_X; reg_b = b7_X; reg_acc = reg_o >> 256; o7_X = reg_o; Enable sign a,b; operation : b +/- a + acc;
"000000100001111000010000001000100001100011111111100010",
--  (2006) addition_subtraction_direct_22
-- NOP 4 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : b + a + acc;
"000000000000000100000000010000011110000100000000000010",
--  (2007) iterative_modular_reduction_0
-- -- In case of size 1
-- reg_a = a0_X; reg_b = 0; reg_acc = 0; Enable sign a,b; operation : b + a + acc;
"000000100001000000000000010000011001100100000000010010",
--  (2008) iterative_modular_reduction_1
-- reg_a = 0; reg_b = prime0; reg_acc = reg_o; reg_s = reg_o_positive; Enable sign a,b; operation : -s*b + a + acc
"000000100001000000000011000111000111100100000000010010",
--  (2009) iterative_modular_reduction_2
-- reg_a = 0; reg_b = prime0; reg_acc = reg_o; reg_s = reg_o_negative; Enable sign a,b; operation : s*b + a + acc
"000000100001000000000001010011000111100100000000010010",
--  (2010) iterative_modular_reduction_3
-- reg_a = 0; reg_b = prime0; reg_acc = reg_o; o0_X = reg_o; reg_s = reg_o_negative; Enable sign a,b; operation : s*b + a + acc
"000000100001000000010001010011000111100100000000010010",
--  (2011) iterative_modular_reduction_4
-- NOP 4 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : b + a + acc;
"000000000000000100000000010000011110000100000000000010",
--  (2012) iterative_modular_reduction_5
-- -- In case of size 2
-- reg_a = a1_X; reg_b = 0; reg_acc = 0; Enable sign a,b; operation : b + a + acc;
"000000100001001000000000010000011001100100000000110010",
--  (2013) iterative_modular_reduction_6
-- reg_a = a0_X; reg_b = prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_positive; operation : -s*b + a + acc
"000000100001001000010011000111010000000100000000010010",
--  (2014) iterative_modular_reduction_7
-- reg_a = a1_X; reg_b = prime1; reg_acc = reg_o >> 256; o1_X = reg_o; Enable sign a,b; operation : -s*b + a + acc
"000000100001001000010011000000100001101000100100110010",
--  (2015) iterative_modular_reduction_8
-- reg_a = o0_X; reg_b = prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc
"000000100001001000010001010011010000000100000000010110",
--  (2016) iterative_modular_reduction_9
-- reg_a = o1_X; reg_b = prime1; reg_acc = reg_o >> 256; o1_X = reg_o; Enable sign a,b operation : s*b + a + acc
"000000100001001000010001010000100001101000100100110110",
--  (2017) iterative_modular_reduction_10
-- reg_a = o0_X; reg_b = prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc
"000000100001001000010001010011010000000100000000010110",
--  (2018) iterative_modular_reduction_11
-- reg_a = o1_X; reg_b = prime1; reg_acc = reg_o >> 256; o1_X = reg_o; Enable sign a,b operation : s*b + a + acc
"000000100001001000010001010000100001101000100100110110",
--  (2019) iterative_modular_reduction_12
-- NOP 4 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : b + a + acc;
"000000000000000100000000010000011110000100000000000010",
--  (2020) iterative_modular_reduction_13
-- -- In case of size 3
-- reg_a = a2_X; reg_b = 0; reg_acc = 0; Enable sign a,b; operation : b + a + acc;
"000000100001010000000000010000011001101101001001010010",
--  (2021) iterative_modular_reduction_14
-- reg_a = a0_X; reg_b = prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_positive; operation : -s*b + a + acc
"000000100001010000010011000111010000000100000000010010",
--  (2022) iterative_modular_reduction_15
-- reg_a = a1_X; reg_b = prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : -s*b + a + acc
"000000100001010000010011000000100000001000100100110010",
--  (2023) iterative_modular_reduction_16
-- reg_a = a2_X; reg_b = prime2; reg_acc = reg_o >> 256; o2_X = reg_o; Enable sign a,b; operation : -s*b + a + acc
"000000100001010000010011000000100001101101001001010010",
--  (2024) iterative_modular_reduction_17
-- reg_a = o0_X; reg_b = prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc
"000000100001010000010001010011010000000100000000010110",
--  (2025) iterative_modular_reduction_18
-- reg_a = o1_X; reg_b = prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : s*b + a + acc
"000000100001010000010001010000100000001000100100110110",
--  (2026) iterative_modular_reduction_19
-- reg_a = o2_X; reg_b = prime2; reg_acc = reg_o >> 256; o2_X = reg_o; Enable sign a,b operation : s*b + a + acc
"000000100001010000010001010000100001101101001001010110",
--  (2027) iterative_modular_reduction_20
-- reg_a = o0_X; reg_b = prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc
"000000100001010000010001010011010000000100000000010110",
--  (2028) iterative_modular_reduction_21
-- reg_a = o1_X; reg_b = prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : s*b + a + acc
"000000100001010000010001010000100000001000100100110110",
--  (2029) iterative_modular_reduction_22
-- reg_a = o2_X; reg_b = prime2; reg_acc = reg_o >> 256; o2_X = reg_o; Enable sign a,b operation : s*b + a + acc
"000000100001010000010001010000100001101101001001010110",
--  (2030) iterative_modular_reduction_23
-- NOP 4 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : b + a + acc;
"000000000000000100000000010000011110000100000000000010",
--  (2031) iterative_modular_reduction_24
-- -- In case of size 4
-- reg_a = a3_X; reg_b = 0; reg_acc = 0; Enable sign a,b; operation : b + a + acc;
"000000100001011000000000010000011001100001101101110010",
--  (2032) iterative_modular_reduction_25
-- reg_a = a0_X; reg_b = prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_positive; operation : -s*b + a + acc
"000000100001011000010011000111010000000100000000010010",
--  (2033) iterative_modular_reduction_26
-- reg_a = a1_X; reg_b = prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : -s*b + a + acc
"000000100001011000010011000000100000001000100100110010",
--  (2034) iterative_modular_reduction_27
-- reg_a = a2_X; reg_b = prime2; reg_acc = reg_o >> 256; o2_X = reg_o; operation : -s*b + a + acc
"000000100001011000010011000000100000001101001001010010",
--  (2035) iterative_modular_reduction_28
-- reg_a = a3_X; reg_b = prime3; reg_acc = reg_o >> 256; o3_X = reg_o; Enable sign a,b; operation : -s*b + a + acc
"000000100001011000010011000000100001100001101101110010",
--  (2036) iterative_modular_reduction_29
-- reg_a = o0_X; reg_b = prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc
"000000100001011000010001010011010000000100000000010110",
--  (2037) iterative_modular_reduction_30
-- reg_a = o1_X; reg_b = prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : s*b + a + acc
"000000100001011000010001010000100000001000100100110110",
--  (2038) iterative_modular_reduction_31
-- reg_a = o2_X; reg_b = prime2; reg_acc = reg_o >> 256; o2_X = reg_o; operation : s*b + a + acc
"000000100001011000010001010000100000001101001001010110",
--  (2039) iterative_modular_reduction_32
-- reg_a = o3_X; reg_b = prime3; reg_acc = reg_o >> 256; o3_X = reg_o; Enable sign a,b; operation : s*b + a + acc
"000000100001011000010001010000100001100001101101110110",
--  (2040) iterative_modular_reduction_33
-- reg_a = o0_X; reg_b = prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc
"000000100001011000010001010011010000000100000000010110",
--  (2041) iterative_modular_reduction_34
-- reg_a = o1_X; reg_b = prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : s*b + a + acc
"000000100001011000010001010000100000001000100100110110",
--  (2042) iterative_modular_reduction_35
-- reg_a = o2_X; reg_b = prime2; reg_acc = reg_o >> 256; o2_X = reg_o; operation : s*b + a + acc
"000000100001011000010001010000100000001101001001010110",
--  (2043) iterative_modular_reduction_36
-- reg_a = o3_X; reg_b = prime3; reg_acc = reg_o >> 256; o3_X = reg_o; Enable sign a,b; operation : s*b + a + acc
"000000100001011000010001010000100001100001101101110110",
--  (2044) iterative_modular_reduction_37
-- NOP 4 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : b + a + acc;
"000000000000000100000000010000011110000100000000000010",
--  (2045) iterative_modular_reduction_38
-- -- In case of size 5
-- reg_a = a4_X; reg_b = 0; reg_acc = 0; Enable sign a,b; operation : b + a + acc;
"000000100001100000000000010000011001110110010010010010",
--  (2046) iterative_modular_reduction_39
-- reg_a = a0_X; reg_b = prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_positive; operation : -s*b + a + acc
"000000100001100000010011000111010000000100000000010010",
--  (2047) iterative_modular_reduction_40
-- reg_a = a1_X; reg_b = prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : -s*b + a + acc
"000000100001100000010011000000100000001000100100110010",
--  (2048) iterative_modular_reduction_41
-- reg_a = a2_X; reg_b = prime2; reg_acc = reg_o >> 256; o2_X = reg_o; operation : -s*b + a + acc
"000000100001100000010011000000100000001101001001010010",
--  (2049) iterative_modular_reduction_42
-- reg_a = a3_X; reg_b = prime3; reg_acc = reg_o >> 256; o3_X = reg_o; operation : -s*b + a + acc
"000000100001100000010011000000100000010001101101110010",
--  (2050) iterative_modular_reduction_43
-- reg_a = a4_X; reg_b = prime4; reg_acc = reg_o >> 256; o4_X = reg_o; Enable sign a,b; operation : -s*b + a + acc
"000000100001100000010011000000100001110110010010010010",
--  (2051) iterative_modular_reduction_44
-- reg_a = o0_X; reg_b = prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc
"000000100001100000010001010011010000000100000000010110",
--  (2052) iterative_modular_reduction_45
-- reg_a = o1_X; reg_b = prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : s*b + a + acc
"000000100001100000010001010000100000001000100100110110",
--  (2053) iterative_modular_reduction_46
-- reg_a = o2_X; reg_b = prime2; reg_acc = reg_o >> 256; o2_X = reg_o; operation : s*b + a + acc
"000000100001100000010001010000100000001101001001010110",
--  (2054) iterative_modular_reduction_47
-- reg_a = o3_X; reg_b = prime3; reg_acc = reg_o >> 256; o3_X = reg_o; operation : s*b + a + acc
"000000100001100000010001010000100000010001101101110110",
--  (2055) iterative_modular_reduction_48
-- reg_a = o4_X; reg_b = prime4; reg_acc = reg_o >> 256; o4_X = reg_o; Enable sign a,b; operation : s*b + a + acc
"000000100001100000010001010000100001110110010010010110",
--  (2056) iterative_modular_reduction_49
-- reg_a = o0_X; reg_b = prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc
"000000100001100000010001010011010000000100000000010110",
--  (2057) iterative_modular_reduction_50
-- reg_a = o1_X; reg_b = prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : s*b + a + acc
"000000100001100000010001010000100000001000100100110110",
--  (2058) iterative_modular_reduction_51
-- reg_a = o2_X; reg_b = prime2; reg_acc = reg_o >> 256; o2_X = reg_o; operation : s*b + a + acc
"000000100001100000010001010000100000001101001001010110",
--  (2059) iterative_modular_reduction_52
-- reg_a = o3_X; reg_b = prime3; reg_acc = reg_o >> 256; o3_X = reg_o; operation : s*b + a + acc
"000000100001100000010001010000100000010001101101110110",
--  (2060) iterative_modular_reduction_53
-- reg_a = o4_X; reg_b = prime4; reg_acc = reg_o >> 256; o4_X = reg_o; Enable sign a,b; operation : s*b + a + acc
"000000100001100000010001010000100001110110010010010110",
--  (2061) iterative_modular_reduction_54
-- NOP 4 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : b + a + acc;
"000000000000000100000000010000011110000100000000000010",
--  (2062) iterative_modular_reduction_55
-- -- In case of size 6
-- reg_a = a5_X; reg_b = 0; reg_acc = 0; Enable sign a,b; operation : b + a + acc;
"000000100001101000000000010000011001111010110110110010",
--  (2063) iterative_modular_reduction_56
-- reg_a = a0_X; reg_b = prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_positive; operation : -s*b + a + acc
"000000100001101000010011000111010000000100000000010010",
--  (2064) iterative_modular_reduction_57
-- reg_a = a1_X; reg_b = prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : -s*b + a + acc
"000000100001101000010011000000100000001000100100110010",
--  (2065) iterative_modular_reduction_58
-- reg_a = a2_X; reg_b = prime2; reg_acc = reg_o >> 256; o2_X = reg_o; operation : -s*b + a + acc
"000000100001101000010011000000100000001101001001010010",
--  (2066) iterative_modular_reduction_59
-- reg_a = a3_X; reg_b = prime3; reg_acc = reg_o >> 256; o3_X = reg_o; operation : -s*b + a + acc
"000000100001101000010011000000100000010001101101110010",
--  (2067) iterative_modular_reduction_60
-- reg_a = a4_X; reg_b = prime4; reg_acc = reg_o >> 256; o4_X = reg_o; operation : -s*b + a + acc
"000000100001101000010011000000100000010110010010010010",
--  (2068) iterative_modular_reduction_61
-- reg_a = a5_X; reg_b = prime5; reg_acc = reg_o >> 256; o5_X = reg_o; Enable sign a,b; operation : -s*b + a + acc
"000000100001101000010011000000100001111010110110110010",
--  (2069) iterative_modular_reduction_62
-- reg_a = o0_X; reg_b = prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc
"000000100001101000010001010011010000000100000000010110",
--  (2070) iterative_modular_reduction_63
-- reg_a = o1_X; reg_b = prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : s*b + a + acc
"000000100001101000010001010000100000001000100100110110",
--  (2071) iterative_modular_reduction_64
-- reg_a = o2_X; reg_b = prime2; reg_acc = reg_o >> 256; o2_X = reg_o; operation : s*b + a + acc
"000000100001101000010001010000100000001101001001010110",
--  (2072) iterative_modular_reduction_65
-- reg_a = o3_X; reg_b = prime3; reg_acc = reg_o >> 256; o3_X = reg_o; operation : s*b + a + acc
"000000100001101000010001010000100000010001101101110110",
--  (2073) iterative_modular_reduction_66
-- reg_a = o4_X; reg_b = prime4; reg_acc = reg_o >> 256; o4_X = reg_o; operation : s*b + a + acc
"000000100001101000010001010000100000010110010010010110",
--  (2074) iterative_modular_reduction_67
-- reg_a = o5_X; reg_b = prime5; reg_acc = reg_o >> 256; o5_X = reg_o; Enable sign a,b; operation : s*b + a + acc
"000000100001101000010001010000100001111010110110110110",
--  (2075) iterative_modular_reduction_68
-- reg_a = o0_X; reg_b = prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc
"000000100001101000010001010011010000000100000000010110",
--  (2076) iterative_modular_reduction_69
-- reg_a = o1_X; reg_b = prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : s*b + a + acc
"000000100001101000010001010000100000001000100100110110",
--  (2077) iterative_modular_reduction_70
-- reg_a = o2_X; reg_b = prime2; reg_acc = reg_o >> 256; o2_X = reg_o; operation : s*b + a + acc
"000000100001101000010001010000100000001101001001010110",
--  (2078) iterative_modular_reduction_71
-- reg_a = o3_X; reg_b = prime3; reg_acc = reg_o >> 256; o3_X = reg_o; operation : s*b + a + acc
"000000100001101000010001010000100000010001101101110110",
--  (2079) iterative_modular_reduction_72
-- reg_a = o4_X; reg_b = prime4; reg_acc = reg_o >> 256; o4_X = reg_o; operation : s*b + a + acc
"000000100001101000010001010000100000010110010010010110",
--  (2080) iterative_modular_reduction_73
-- reg_a = o5_X; reg_b = prime5; reg_acc = reg_o >> 256; o5_X = reg_o; Enable sign a,b; operation : s*b + a + acc
"000000100001101000010001010000100001111010110110110110",
--  (2081) iterative_modular_reduction_74
-- NOP 4 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : b + a + acc;
"000000000000000100000000010000011110000100000000000010",
--  (2082) iterative_modular_reduction_75
-- -- In case of size 7
-- reg_a = a6_X; reg_b = 0; reg_acc = 0; Enable sign a,b; operation : b + a + acc;
"000000100001110000000000010000011001111111011011010010",
--  (2083) iterative_modular_reduction_76
-- reg_a = a0_X; reg_b = prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_positive; operation : -s*b + a + acc
"000000100001110000010011000111010000000100000000010010",
--  (2084) iterative_modular_reduction_77
-- reg_a = a1_X; reg_b = prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : -s*b + a + acc
"000000100001110000010011000000100000001000100100110010",
--  (2085) iterative_modular_reduction_78
-- reg_a = a2_X; reg_b = prime2; reg_acc = reg_o >> 256; o2_X = reg_o; operation : -s*b + a + acc
"000000100001110000010011000000100000001101001001010010",
--  (2086) iterative_modular_reduction_79
-- reg_a = a3_X; reg_b = prime3; reg_acc = reg_o >> 256; o3_X = reg_o; operation : -s*b + a + acc
"000000100001110000010011000000100000010001101101110010",
--  (2087) iterative_modular_reduction_80
-- reg_a = a4_X; reg_b = prime4; reg_acc = reg_o >> 256; o4_X = reg_o; operation : -s*b + a + acc
"000000100001110000010011000000100000010110010010010010",
--  (2088) iterative_modular_reduction_81
-- reg_a = a5_X; reg_b = prime5; reg_acc = reg_o >> 256; o5_X = reg_o; operation : -s*b + a + acc
"000000100001110000010011000000100000011010110110110010",
--  (2089) iterative_modular_reduction_82
-- reg_a = a6_X; reg_b = prime6; reg_acc = reg_o >> 256; o6_X = reg_o; Enable sign a,b; operation : -s*b + a + acc
"000000100001110000010011000000100001111111011011010010",
--  (2090) iterative_modular_reduction_83
-- reg_a = o0_X; reg_b = prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc
"000000100001110000010001010011010000000100000000010110",
--  (2091) iterative_modular_reduction_84
-- reg_a = o1_X; reg_b = prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : s*b + a + acc
"000000100001110000010001010000100000001000100100110110",
--  (2092) iterative_modular_reduction_85
-- reg_a = o2_X; reg_b = prime2; reg_acc = reg_o >> 256; o2_X = reg_o; operation : s*b + a + acc
"000000100001110000010001010000100000001101001001010110",
--  (2093) iterative_modular_reduction_86
-- reg_a = o3_X; reg_b = prime3; reg_acc = reg_o >> 256; o3_X = reg_o; operation : s*b + a + acc
"000000100001110000010001010000100000010001101101110110",
--  (2094) iterative_modular_reduction_87
-- reg_a = o4_X; reg_b = prime4; reg_acc = reg_o >> 256; o4_X = reg_o; operation : s*b + a + acc
"000000100001110000010001010000100000010110010010010110",
--  (2095) iterative_modular_reduction_88
-- reg_a = o5_X; reg_b = prime5; reg_acc = reg_o >> 256; o5_X = reg_o; operation : s*b + a + acc
"000000100001110000010001010000100000011010110110110110",
--  (2096) iterative_modular_reduction_89
-- reg_a = o6_X; reg_b = prime6; reg_acc = reg_o >> 256; o6_X = reg_o; Enable sign a,b; operation : s*b + a + acc
"000000100001110000010001010000100001111111011011010110",
--  (2097) iterative_modular_reduction_90
-- reg_a = o0_X; reg_b = prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc
"000000100001110000010001010011010000000100000000010110",
--  (2098) iterative_modular_reduction_91
-- reg_a = o1_X; reg_b = prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : s*b + a + acc
"000000100001110000010001010000100000001000100100110110",
--  (2099) iterative_modular_reduction_92
-- reg_a = o2_X; reg_b = prime2; reg_acc = reg_o >> 256; o2_X = reg_o; operation : s*b + a + acc
"000000100001110000010001010000100000001101001001010110",
--  (2100) iterative_modular_reduction_93
-- reg_a = o3_X; reg_b = prime3; reg_acc = reg_o >> 256; o3_X = reg_o; operation : s*b + a + acc
"000000100001110000010001010000100000010001101101110110",
--  (2101) iterative_modular_reduction_94
-- reg_a = o4_X; reg_b = prime4; reg_acc = reg_o >> 256; o4_X = reg_o; operation : s*b + a + acc
"000000100001110000010001010000100000010110010010010110",
--  (2102) iterative_modular_reduction_95
-- reg_a = o5_X; reg_b = prime5; reg_acc = reg_o >> 256; o5_X = reg_o; operation : s*b + a + acc
"000000100001110000010001010000100000011010110110110110",
--  (2103) iterative_modular_reduction_96
-- reg_a = o6_X; reg_b = prime6; reg_acc = reg_o >> 256; o6_X = reg_o; Enable sign a,b; operation : s*b + a + acc
"000000100001110000010001010000100001111111011011010110",
--  (2104) iterative_modular_reduction_97
-- NOP 4 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : b + a + acc;
"000000000000000100000000010000011110000100000000000010",
--  (2105) iterative_modular_reduction_98
-- -- In case of size 8
-- reg_a = a7_X; reg_b = 0; reg_acc = 0; Enable sign a,b; operation : b + a + acc;
"000000100001111000000000010000011001100011111111110010",
--  (2106) iterative_modular_reduction_99
-- reg_a = a0_X; reg_b = prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_positive; operation : -s*b + a + acc
"000000100001111000010011000111010000000100000000010010",
--  (2107) iterative_modular_reduction_100
-- reg_a = a1_X; reg_b = prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : -s*b + a + acc
"000000100001111000010011000000100000001000100100110010",
--  (2108) iterative_modular_reduction_101
-- reg_a = a2_X; reg_b = prime2; reg_acc = reg_o >> 256; o2_X = reg_o; operation : -s*b + a + acc
"000000100001111000010011000000100000001101001001010010",
--  (2109) iterative_modular_reduction_102
-- reg_a = a3_X; reg_b = prime3; reg_acc = reg_o >> 256; o3_X = reg_o; operation : -s*b + a + acc
"000000100001111000010011000000100000010001101101110010",
--  (2110) iterative_modular_reduction_103
-- reg_a = a4_X; reg_b = prime4; reg_acc = reg_o >> 256; o4_X = reg_o; operation : -s*b + a + acc
"000000100001111000010011000000100000010110010010010010",
--  (2111) iterative_modular_reduction_104
-- reg_a = a5_X; reg_b = prime5; reg_acc = reg_o >> 256; o5_X = reg_o; operation : -s*b + a + acc
"000000100001111000010011000000100000011010110110110010",
--  (2112) iterative_modular_reduction_105
-- reg_a = a6_X; reg_b = prime6; reg_acc = reg_o >> 256; o6_X = reg_o; operation : -s*b + a + acc
"000000100001111000010011000000100000011111011011010010",
--  (2113) iterative_modular_reduction_106
-- reg_a = a7_X; reg_b = prime7; reg_acc = reg_o >> 256; o7_X = reg_o; Enable sign a,b; operation : -s*b + a + acc
"000000100001111000010011000000100001100011111111110010",
--  (2114) iterative_modular_reduction_107
-- reg_a = o0_X; reg_b = prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc
"000000100001111000010001010011010000000100000000010110",
--  (2115) iterative_modular_reduction_108
-- reg_a = o1_X; reg_b = prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : s*b + a + acc
"000000100001111000010001010000100000001000100100110110",
--  (2116) iterative_modular_reduction_109
-- reg_a = o2_X; reg_b = prime2; reg_acc = reg_o >> 256; o2_X = reg_o; operation : s*b + a + acc
"000000100001111000010001010000100000001101001001010110",
--  (2117) iterative_modular_reduction_110
-- reg_a = o3_X; reg_b = prime3; reg_acc = reg_o >> 256; o3_X = reg_o; operation : s*b + a + acc
"000000100001111000010001010000100000010001101101110110",
--  (2118) iterative_modular_reduction_111
-- reg_a = o4_X; reg_b = prime4; reg_acc = reg_o >> 256; o4_X = reg_o; operation : s*b + a + acc
"000000100001111000010001010000100000010110010010010110",
--  (2119) iterative_modular_reduction_112
-- reg_a = o5_X; reg_b = prime5; reg_acc = reg_o >> 256; o5_X = reg_o; operation : s*b + a + acc
"000000100001111000010001010000100000011010110110110110",
--  (2120) iterative_modular_reduction_113
-- reg_a = o6_X; reg_b = prime6; reg_acc = reg_o >> 256; o6_X = reg_o; operation : s*b + a + acc
"000000100001111000010001010000100000011111011011010110",
--  (2121) iterative_modular_reduction_114
-- reg_a = o7_X; reg_b = prime7; reg_acc = reg_o >> 256; o7_X = reg_o; Enable sign a,b; operation : s*b + a + acc
"000000100001111000010001010000100001100011111111110110",
--  (2122) iterative_modular_reduction_115
-- reg_a = o0_X; reg_b = prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc
"000000100001111000010001010011010000000100000000010110",
--  (2123) iterative_modular_reduction_116
-- reg_a = o1_X; reg_b = prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : s*b + a + acc
"000000100001111000010001010000100000001000100100110110",
--  (2124) iterative_modular_reduction_117
-- reg_a = o2_X; reg_b = prime2; reg_acc = reg_o >> 256; o2_X = reg_o; operation : s*b + a + acc
"000000100001111000010001010000100000001101001001010110",
--  (2125) iterative_modular_reduction_118
-- reg_a = o3_X; reg_b = prime3; reg_acc = reg_o >> 256; o3_X = reg_o; operation : s*b + a + acc
"000000100001111000010001010000100000010001101101110110",
--  (2126) iterative_modular_reduction_119
-- reg_a = o4_X; reg_b = prime4; reg_acc = reg_o >> 256; o4_X = reg_o; operation : s*b + a + acc
"000000100001111000010001010000100000010110010010010110",
--  (2127) iterative_modular_reduction_120
-- reg_a = o5_X; reg_b = prime5; reg_acc = reg_o >> 256; o5_X = reg_o; operation : s*b + a + acc
"000000100001111000010001010000100000011010110110110110",
--  (2128) iterative_modular_reduction_121
-- reg_a = o6_X; reg_b = prime6; reg_acc = reg_o >> 256; o6_X = reg_o; operation : s*b + a + acc
"000000100001111000010001010000100000011111011011010110",
--  (2129) iterative_modular_reduction_122
-- reg_a = o7_X; reg_b = prime7; reg_acc = reg_o >> 256; o7_X = reg_o; Enable sign a,b; operation : s*b + a + acc
"000000100001111000010001010000100001100011111111110110",
--  (2130) iterative_modular_reduction_123
-- NOP 4 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : b + a + acc;
"000000000000000100000000010000011110000100000000000010",
--  (2131) addition_subtraction_with_reduction_0
-- Operands size 1
-- reg_a = a0_X; reg_b = b0_X; reg_acc = 0; o0_X = reg_o; Enable sign a,b; operation : b +/- a + acc;
"000000100001000000010000011000010001100100000000000010",
--  (2132) addition_subtraction_with_reduction_1
-- reg_a = 0; reg_b = 2prime0; reg_acc = reg_o; reg_s = reg_o_positive; o0_X = reg_o; Enable sign a,b; operation : -s*b + a + acc;
"000000100001000000010011000111000111100100000000001010",
--  (2133) addition_subtraction_with_reduction_2
-- reg_a = 0; reg_b = 2prime0; reg_acc = reg_o; reg_s = reg_o_negative; o0_X = reg_o; Enable sign a,b; operation : s*b + a + acc;
"000000100001000000010001010011000111100100000000001010",
--  (2134) addition_subtraction_with_reduction_3
-- reg_a = 0; reg_b = 2prime0; reg_acc = reg_o; reg_s = reg_o_negative; o0_X = reg_o; Enable sign a,b; operation : s*b + a + acc;
"000000100001000000010001010011000111100100000000001010",
--  (2135) addition_subtraction_with_reduction_4
-- NOP 4 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : b + a + acc;
"000000000000000100000000010000011110000100000000000010",
--  (2136) addition_subtraction_with_reduction_5
-- -- In case of sizes 2, 3, 4, 5, 6, 7, 8
-- reg_a = a0_X; reg_b = b0_X; reg_acc = 0; o0_X = reg_o; operation : b +/- a + acc;
"000100100001001000010000001000010000000100000000000010",
--  (2137) addition_subtraction_with_reduction_6
-- -- In case of size 2
-- reg_a = a1_X; reg_b = b1_X; reg_acc = reg_o >> 256; o1_X = reg_o; Enable sign a, b; operation : b +/- a + acc;
"000000100001001000010000001000100001101000100100100010",
--  (2138) addition_subtraction_with_reduction_7
-- reg_a = o0_X; reg_b = 2prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_positive; operation : -s*b + a + acc;
"000000100001001000010011000111010000000100000000001110",
--  (2139) addition_subtraction_with_reduction_8
-- reg_a = o1_X; reg_b = 2prime1; reg_acc = reg_o >> 256; o1_X = reg_o; Enable sign a,b; operation : -s*b + a + acc;
"000000100001001000010011000000100001101000100100101110",
--  (2140) addition_subtraction_with_reduction_9
-- reg_a = o0_X; reg_b = 2prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc;
"000000100001001000010001010011010000000100000000001110",
--  (2141) addition_subtraction_with_reduction_10
-- reg_a = o1_X; reg_b = 2prime1; reg_acc = reg_o >> 256; o1_X = reg_o; Enable sign a,b; operation : s*b + a + acc;
"000000100001001000010001010000100001101000100100101110",
--  (2142) addition_subtraction_with_reduction_11
-- reg_a = o0_X; reg_b = 2prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc;
"000000100001001000010001010011010000000100000000001110",
--  (2143) addition_subtraction_with_reduction_12
-- reg_a = o1_X; reg_b = 2prime1; reg_acc = reg_o >> 256; o1_X = reg_o; Enable sign a,b; operation : s*b + a + acc;
"000000100001001000010001010000100001101000100100101110",
--  (2144) addition_subtraction_with_reduction_13
-- NOP 4 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : b + a + acc;
"000000000000000100000000010000011110000100000000000010",
--  (2145) addition_subtraction_with_reduction_14
-- -- In case of sizes 3, 4, 5, 6, 7, 8
-- reg_a = a1_X; reg_b = b1_X; reg_acc = reg_o >> 256; o1_X = reg_o; operation : b +/- a + acc;
"000110000001010000010000001000100000001000100100100010",
--  (2146) addition_subtraction_with_reduction_15
-- -- In case of size 3
-- reg_a = a2_X; reg_b = b2_X; reg_acc = reg_o >> 256; o2_X = reg_o; Enable sign a, b; operation : b +/- a + acc;
"000000100001010000010000001000100001100101001001000010",
--  (2147) addition_subtraction_with_reduction_16
-- reg_a = o0_X; reg_b = 2prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_positive; operation : -s*b + a + acc;
"000000100001010000010011000111010000000100000000001110",
--  (2148) addition_subtraction_with_reduction_17
-- reg_a = o1_X; reg_b = 2prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : -s*b + a + acc;
"000000100001010000010011000000100000001000100100101110",
--  (2149) addition_subtraction_with_reduction_18
-- reg_a = o2_X; reg_b = 2prime2; reg_acc = reg_o >> 256; o2_X = reg_o; Enable sign a,b; operation : -s*b + a + acc;
"000000100001010000010011000000100001101101001001001110",
--  (2150) addition_subtraction_with_reduction_19
-- reg_a = o0_X; reg_b = 2prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc;
"000000100001010000010001010011010000000100000000001110",
--  (2151) addition_subtraction_with_reduction_20
-- reg_a = o1_X; reg_b = 2prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : s*b + a + acc;
"000000100001010000010001010000100000001000100100101110",
--  (2152) addition_subtraction_with_reduction_21
-- reg_a = o2_X; reg_b = 2prime2; reg_acc = reg_o >> 256; o2_X = reg_o; Enable sign a,b; operation : s*b + a + acc;
"000000100001010000010001010000100001101101001001001110",
--  (2153) addition_subtraction_with_reduction_22
-- reg_a = o0_X; reg_b = 2prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc;
"000000100001010000010001010011010000000100000000001110",
--  (2154) addition_subtraction_with_reduction_23
-- reg_a = o1_X; reg_b = 2prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : s*b + a + acc;
"000000100001010000010001010000100000001000100100101110",
--  (2155) addition_subtraction_with_reduction_24
-- reg_a = o2_X; reg_b = 2prime2; reg_acc = reg_o >> 256; o2_X = reg_o; Enable sign a,b; operation : s*b + a + acc;
"000000100001010000010001010000100001101101001001001110",
--  (2156) addition_subtraction_with_reduction_25
-- NOP 4 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : b + a + acc;
"000000000000000100000000010000011110000100000000000010",
--  (2157) addition_subtraction_with_reduction_26
-- -- In case of size 4, 5, 6, 7, 8
-- reg_a = a2_X; reg_b = b2_X; reg_acc = reg_o >> 256; o2_X = reg_o; operation : b +/- a + acc;
"000111100001011000010000001000100000000101001001000010",
--  (2158) addition_subtraction_with_reduction_27
-- -- In case of size 4
-- reg_a = a3_X; reg_b = b3_X; reg_acc = reg_o >> 256; o3_X = reg_o; Enable sign a, b; operation : b +/- a + acc;
"000000100001011000010000001000100001110001101101100010",
--  (2159) addition_subtraction_with_reduction_28
-- reg_a = o0_X; reg_b = 2prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_positive; operation : -s*b + a + acc;
"000000100001011000010011000111010000000100000000001110",
--  (2160) addition_subtraction_with_reduction_29
-- reg_a = o1_X; reg_b = 2prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : -s*b + a + acc;
"000000100001011000010011000000100000001000100100101110",
--  (2161) addition_subtraction_with_reduction_30
-- reg_a = o2_X; reg_b = 2prime2; reg_acc = reg_o >> 256; o2_X = reg_o; operation : -s*b + a + acc;
"000000100001011000010011000000100000001101001001001110",
--  (2162) addition_subtraction_with_reduction_31
-- reg_a = o3_X; reg_b = 2prime3; reg_acc = reg_o >> 256; o3_X = reg_o; Enable sign a,b; operation : -s*b + a + acc;
"000000100001011000010011000000100001100001101101101110",
--  (2163) addition_subtraction_with_reduction_32
-- reg_a = o0_X; reg_b = 2prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc;
"000000100001011000010001010011010000000100000000001110",
--  (2164) addition_subtraction_with_reduction_33
-- reg_a = o1_X; reg_b = 2prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : s*b + a + acc;
"000000100001011000010001010000100000001000100100101110",
--  (2165) addition_subtraction_with_reduction_34
-- reg_a = o2_X; reg_b = 2prime2; reg_acc = reg_o >> 256; o2_X = reg_o; operation : s*b + a + acc;
"000000100001011000010001010000100000001101001001001110",
--  (2166) addition_subtraction_with_reduction_35
-- reg_a = o3_X; reg_b = 2prime3; reg_acc = reg_o >> 256; o3_X = reg_o; Enable sign a,b; operation : s*b + a + acc;
"000000100001011000010001010000100001100001101101101110",
--  (2167) addition_subtraction_with_reduction_36
-- reg_a = o0_X; reg_b = 2prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc;
"000000100001011000010001010011010000000100000000001110",
--  (2168) addition_subtraction_with_reduction_37
-- reg_a = o1_X; reg_b = 2prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : s*b + a + acc;
"000000100001011000010001010000100000001000100100101110",
--  (2169) addition_subtraction_with_reduction_38
-- reg_a = o2_X; reg_b = 2prime2; reg_acc = reg_o >> 256; o2_X = reg_o; operation : s*b + a + acc;
"000000100001011000010001010000100000001101001001001110",
--  (2170) addition_subtraction_with_reduction_39
-- reg_a = o3_X; reg_b = 2prime3; reg_acc = reg_o >> 256; o3_X = reg_o; Enable sign a,b; operation : s*b + a + acc;
"000000100001011000010001010000100001110001101101101110",
--  (2171) addition_subtraction_with_reduction_40
-- NOP 4 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : b + a + acc;
"000000000000000100000000010000011110000100000000000010",
--  (2172) addition_subtraction_with_reduction_41
-- -- In case of size 5, 6, 7, 8
-- reg_a = a3_X; reg_b = b3_X; reg_acc = reg_o >> 256; o3_X = reg_o; operation : b +/- a + acc;
"001001000001100000010000001000100000010001101101100010",
--  (2173) addition_subtraction_with_reduction_42
-- -- In case of size 5
-- reg_a = a4_X; reg_b = b4_X; reg_acc = reg_o >> 256; o4_X = reg_o; Enable sign a, b; operation : b +/- a + acc;
"000000100001100000010000001000100001110110010010000010",
--  (2174) addition_subtraction_with_reduction_43
-- reg_a = o0_X; reg_b = 2prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_positive; operation : -s*b + a + acc;
"000000100001100000010011000111010000000100000000001110",
--  (2175) addition_subtraction_with_reduction_44
-- reg_a = o1_X; reg_b = 2prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : -s*b + a + acc;
"000000100001100000010011000000100000001000100100101110",
--  (2176) addition_subtraction_with_reduction_45
-- reg_a = o2_X; reg_b = 2prime2; reg_acc = reg_o >> 256; o2_X = reg_o; operation : -s*b + a + acc;
"000000100001100000010011000000100000001101001001001110",
--  (2177) addition_subtraction_with_reduction_46
-- reg_a = o3_X; reg_b = 2prime3; reg_acc = reg_o >> 256; o3_X = reg_o; operation : -s*b + a + acc;
"000000100001100000010011000000100000010001101101101110",
--  (2178) addition_subtraction_with_reduction_47
-- reg_a = o4_X; reg_b = 2prime4; reg_acc = reg_o >> 256; o4_X = reg_o; Enable sign a,b; operation : -s*b + a + acc;
"000000100001100000010011000000100001110110010010001110",
--  (2179) addition_subtraction_with_reduction_48
-- reg_a = o0_X; reg_b = 2prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc;
"000000100001100000010001010011010000000100000000001110",
--  (2180) addition_subtraction_with_reduction_49
-- reg_a = o1_X; reg_b = 2prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : s*b + a + acc;
"000000100001100000010001010000100000001000100100101110",
--  (2181) addition_subtraction_with_reduction_50
-- reg_a = o2_X; reg_b = 2prime2; reg_acc = reg_o >> 256; o2_X = reg_o; operation : s*b + a + acc;
"000000100001100000010001010000100000001101001001001110",
--  (2182) addition_subtraction_with_reduction_51
-- reg_a = o3_X; reg_b = 2prime3; reg_acc = reg_o >> 256; o3_X = reg_o; operation : s*b + a + acc;
"000000100001100000010001010000100000010001101101101110",
--  (2183) addition_subtraction_with_reduction_52
-- reg_a = o4_X; reg_b = 2prime4; reg_acc = reg_o >> 256; o4_X = reg_o; Enable sign a,b; operation : s*b + a + acc;
"000000100001100000010001010000100001110110010010001110",
--  (2184) addition_subtraction_with_reduction_53
-- reg_a = o0_X; reg_b = 2prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc;
"000000100001100000010001010011010000000100000000001110",
--  (2185) addition_subtraction_with_reduction_54
-- reg_a = o1_X; reg_b = 2prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : s*b + a + acc;
"000000100001100000010001010000100000001000100100101110",
--  (2186) addition_subtraction_with_reduction_55
-- reg_a = o2_X; reg_b = 2prime2; reg_acc = reg_o >> 256; o2_X = reg_o; operation : s*b + a + acc;
"000000100001100000010001010000100000001101001001001110",
--  (2187) addition_subtraction_with_reduction_56
-- reg_a = o3_X; reg_b = 2prime3; reg_acc = reg_o >> 256; o3_X = reg_o; operation : s*b + a + acc;
"000000100001100000010001010000100000010001101101101110",
--  (2188) addition_subtraction_with_reduction_57
-- reg_a = o4_X; reg_b = 2prime4; reg_acc = reg_o >> 256; o4_X = reg_o; Enable sign a,b; operation : s*b + a + acc;
"000000100001100000010001010000100001110110010010001110",
--  (2189) addition_subtraction_with_reduction_58
-- NOP 4 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : b + a + acc;
"000000000000000100000000010000011110000100000000000010",
--  (2190) addition_subtraction_with_reduction_59
-- -- In case of size 6, 7, 8
-- reg_a = a4_X; reg_b = b4_X; reg_acc = reg_o >> 256; o4_X = reg_o; operation : b +/- a + acc;
"001010100001101000010000001000100000010110010010000010",
--  (2191) addition_subtraction_with_reduction_60
-- -- In case of size 6
-- reg_a = a5_X; reg_b = b5_X; reg_acc = reg_o >> 256; o5_X = reg_o; Enable sign a, b; operation : b +/- a + acc;
"000000100001101000010000001000100001111010110110100010",
--  (2192) addition_subtraction_with_reduction_61
-- reg_a = o0_X; reg_b = 2prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_positive; operation : -s*b + a + acc;
"000000100001101000010011000111010000000100000000001110",
--  (2193) addition_subtraction_with_reduction_62
-- reg_a = o1_X; reg_b = 2prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : -s*b + a + acc;
"000000100001101000010011000000100000001000100100101110",
--  (2194) addition_subtraction_with_reduction_63
-- reg_a = o2_X; reg_b = 2prime2; reg_acc = reg_o >> 256; o2_X = reg_o; operation : -s*b + a + acc;
"000000100001101000010011000000100000001101001001001110",
--  (2195) addition_subtraction_with_reduction_64
-- reg_a = o3_X; reg_b = 2prime3; reg_acc = reg_o >> 256; o3_X = reg_o; operation : -s*b + a + acc;
"000000100001101000010011000000100000010001101101101110",
--  (2196) addition_subtraction_with_reduction_65
-- reg_a = o4_X; reg_b = 2prime4; reg_acc = reg_o >> 256; o4_X = reg_o; operation : -s*b + a + acc;
"000000100001101000010011000000100000010110010010001110",
--  (2197) addition_subtraction_with_reduction_66
-- reg_a = o5_X; reg_b = 2prime5; reg_acc = reg_o >> 256; o5_X = reg_o; Enable sign a,b; operation : -s*b + a + acc;
"000000100001101000010011000000100001111010110110101110",
--  (2198) addition_subtraction_with_reduction_67
-- reg_a = o0_X; reg_b = 2prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc;
"000000100001101000010001010011010000000100000000001110",
--  (2199) addition_subtraction_with_reduction_68
-- reg_a = o1_X; reg_b = 2prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : s*b + a + acc;
"000000100001101000010001010000100000001000100100101110",
--  (2200) addition_subtraction_with_reduction_69
-- reg_a = o2_X; reg_b = 2prime2; reg_acc = reg_o >> 256; o2_X = reg_o; operation : s*b + a + acc;
"000000100001101000010001010000100000001101001001001110",
--  (2201) addition_subtraction_with_reduction_70
-- reg_a = o3_X; reg_b = 2prime3; reg_acc = reg_o >> 256; o3_X = reg_o; operation : s*b + a + acc;
"000000100001101000010001010000100000010001101101101110",
--  (2202) addition_subtraction_with_reduction_71
-- reg_a = o4_X; reg_b = 2prime4; reg_acc = reg_o >> 256; o4_X = reg_o; operation : s*b + a + acc;
"000000100001101000010001010000100000010110010010001110",
--  (2203) addition_subtraction_with_reduction_72
-- reg_a = o5_X; reg_b = 2prime5; reg_acc = reg_o >> 256; o5_X = reg_o; Enable sign a,b; operation : s*b + a + acc;
"000000100001101000010001010000100001111010110110101110",
--  (2204) addition_subtraction_with_reduction_73
-- reg_a = o0_X; reg_b = 2prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc;
"000000100001101000010001010011010000000100000000001110",
--  (2205) addition_subtraction_with_reduction_74
-- reg_a = o1_X; reg_b = 2prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : s*b + a + acc;
"000000100001101000010001010000100000001000100100101110",
--  (2206) addition_subtraction_with_reduction_75
-- reg_a = o2_X; reg_b = 2prime2; reg_acc = reg_o >> 256; o2_X = reg_o; operation : s*b + a + acc;
"000000100001101000010001010000100000001101001001001110",
--  (2207) addition_subtraction_with_reduction_76
-- reg_a = o3_X; reg_b = 2prime3; reg_acc = reg_o >> 256; o3_X = reg_o; operation : s*b + a + acc;
"000000100001101000010001010000100000010001101101101110",
--  (2208) addition_subtraction_with_reduction_77
-- reg_a = o4_X; reg_b = 2prime4; reg_acc = reg_o >> 256; o4_X = reg_o; operation : s*b + a + acc;
"000000100001101000010001010000100000010110010010001110",
--  (2209) addition_subtraction_with_reduction_78
-- reg_a = o5_X; reg_b = 2prime5; reg_acc = reg_o >> 256; o5_X = reg_o; Enable sign a,b; operation : s*b + a + acc;
"000000100001101000010001010000100001111010110110101110",
--  (2210) addition_subtraction_with_reduction_79
-- NOP 4 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : b + a + acc;
"000000000000000100000000010000011110000100000000000010",
--  (2211) addition_subtraction_with_reduction_80
-- -- In case of size 7, 8
-- reg_a = a5_X; reg_b = b5_X; reg_acc = reg_o >> 256; o5_X = reg_o; operation : b +/- a + acc;
"001100000001110000010000001000100000011010110110100010",
--  (2212) addition_subtraction_with_reduction_81
-- -- In case of size 7
-- reg_a = a6_X; reg_b = b6_X; reg_acc = reg_o >> 256; o6_X = reg_o; Enable sign a, b; operation : b +/- a + acc;
"000000100001110000010000001000100001111111011011000010",
--  (2213) addition_subtraction_with_reduction_82
-- reg_a = o0_X; reg_b = 2prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_positive; operation : -s*b + a + acc;
"000000100001110000010011000111010000000100000000001110",
--  (2214) addition_subtraction_with_reduction_83
-- reg_a = o1_X; reg_b = 2prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : -s*b + a + acc;
"000000100001110000010011000000100000001000100100101110",
--  (2215) addition_subtraction_with_reduction_84
-- reg_a = o2_X; reg_b = 2prime2; reg_acc = reg_o >> 256; o2_X = reg_o; operation : -s*b + a + acc;
"000000100001110000010011000000100000001101001001001110",
--  (2216) addition_subtraction_with_reduction_85
-- reg_a = o3_X; reg_b = 2prime3; reg_acc = reg_o >> 256; o3_X = reg_o; operation : -s*b + a + acc;
"000000100001110000010011000000100000010001101101101110",
--  (2217) addition_subtraction_with_reduction_86
-- reg_a = o4_X; reg_b = 2prime4; reg_acc = reg_o >> 256; o4_X = reg_o; operation : -s*b + a + acc;
"000000100001110000010011000000100000010110010010001110",
--  (2218) addition_subtraction_with_reduction_87
-- reg_a = o5_X; reg_b = 2prime5; reg_acc = reg_o >> 256; o5_X = reg_o; operation : -s*b + a + acc;
"000000100001110000010011000000100000011010110110101110",
--  (2219) addition_subtraction_with_reduction_88
-- reg_a = o6_X; reg_b = 2prime6; reg_acc = reg_o >> 256; o6_X = reg_o; Enable sign a,b; operation : -s*b + a + acc;
"000000100001110000010011000000100001111111011011001110",
--  (2220) addition_subtraction_with_reduction_89
-- reg_a = o0_X; reg_b = 2prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc;
"000000100001110000010001010011010000000100000000001110",
--  (2221) addition_subtraction_with_reduction_90
-- reg_a = o1_X; reg_b = 2prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : s*b + a + acc;
"000000100001110000010001010000100000001000100100101110",
--  (2222) addition_subtraction_with_reduction_91
-- reg_a = o2_X; reg_b = 2prime2; reg_acc = reg_o >> 256; o2_X = reg_o; operation : s*b + a + acc;
"000000100001110000010001010000100000001101001001001110",
--  (2223) addition_subtraction_with_reduction_92
-- reg_a = o3_X; reg_b = 2prime3; reg_acc = reg_o >> 256; o3_X = reg_o; operation : s*b + a + acc;
"000000100001110000010001010000100000010001101101101110",
--  (2224) addition_subtraction_with_reduction_93
-- reg_a = o4_X; reg_b = 2prime4; reg_acc = reg_o >> 256; o4_X = reg_o; operation : s*b + a + acc;
"000000100001110000010001010000100000010110010010001110",
--  (2225) addition_subtraction_with_reduction_94
-- reg_a = o5_X; reg_b = 2prime5; reg_acc = reg_o >> 256; o5_X = reg_o; operation : s*b + a + acc;
"000000100001110000010001010000100000011010110110101110",
--  (2226) addition_subtraction_with_reduction_95
-- reg_a = o6_X; reg_b = 2prime6; reg_acc = reg_o >> 256; o6_X = reg_o; Enable sign a,b; operation : s*b + a + acc;
"000000100001110000010001010000100001111111011011001110",
--  (2227) addition_subtraction_with_reduction_96
-- reg_a = o0_X; reg_b = 2prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc;
"000000100001110000010001010011010000000100000000001110",
--  (2228) addition_subtraction_with_reduction_97
-- reg_a = o1_X; reg_b = 2prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : s*b + a + acc;
"000000100001110000010001010000100000001000100100101110",
--  (2229) addition_subtraction_with_reduction_98
-- reg_a = o2_X; reg_b = 2prime2; reg_acc = reg_o >> 256; o2_X = reg_o; operation : s*b + a + acc;
"000000100001110000010001010000100000001101001001001110",
--  (2230) addition_subtraction_with_reduction_99
-- reg_a = o3_X; reg_b = 2prime3; reg_acc = reg_o >> 256; o3_X = reg_o; operation : s*b + a + acc;
"000000100001110000010001010000100000010001101101101110",
--  (2231) addition_subtraction_with_reduction_100
-- reg_a = o4_X; reg_b = 2prime4; reg_acc = reg_o >> 256; o4_X = reg_o; operation : s*b + a + acc;
"000000100001110000010001010000100000010110010010001110",
--  (2232) addition_subtraction_with_reduction_101
-- reg_a = o5_X; reg_b = 2prime5; reg_acc = reg_o >> 256; o5_X = reg_o; operation : s*b + a + acc;
"000000100001110000010001010000100000011010110110101110",
--  (2233) addition_subtraction_with_reduction_102
-- reg_a = o6_X; reg_b = 2prime6; reg_acc = reg_o >> 256; o6_X = reg_o; Enable sign a,b; operation : s*b + a + acc;
"000000100001110000010001010000100001111111011011001110",
--  (2234) addition_subtraction_with_reduction_103
-- NOP 4 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : b + a + acc;
"000000000000000100000000010000011110000100000000000010",
--  (2235) addition_subtraction_with_reduction_104
-- -- In case of size 8
-- reg_a = a6_X; reg_b = b6_X; reg_acc = reg_o >> 256; o6_X = reg_o; operation : b +/- a + acc;
"000000100001111000010000001000100000011111011011000010",
--  (2236) addition_subtraction_with_reduction_105
-- reg_a = a7_X; reg_b = b7_X; reg_acc = reg_o >> 256; o7_X = reg_o; Enable sign a,b; operation : b +/- a + acc;
"000000100001111000010000001000100001100011111111100010",
--  (2237) addition_subtraction_with_reduction_106
-- reg_a = o0_X; reg_b = 2prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_positive; operation : -s*b + a + acc;
"000000100001111000010011000111010000000100000000001110",
--  (2238) addition_subtraction_with_reduction_107
-- reg_a = o1_X; reg_b = 2prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : -s*b + a + acc;
"000000100001111000010011000000100000001000100100101110",
--  (2239) addition_subtraction_with_reduction_108
-- reg_a = o2_X; reg_b = 2prime2; reg_acc = reg_o >> 256; o2_X = reg_o; operation : -s*b + a + acc;
"000000100001111000010011000000100000001101001001001110",
--  (2240) addition_subtraction_with_reduction_109
-- reg_a = o3_X; reg_b = 2prime3; reg_acc = reg_o >> 256; o3_X = reg_o; operation : -s*b + a + acc;
"000000100001111000010011000000100000010001101101101110",
--  (2241) addition_subtraction_with_reduction_110
-- reg_a = o4_X; reg_b = 2prime4; reg_acc = reg_o >> 256; o4_X = reg_o; operation : -s*b + a + acc;
"000000100001111000010011000000100000010110010010001110",
--  (2242) addition_subtraction_with_reduction_111
-- reg_a = o5_X; reg_b = 2prime5; reg_acc = reg_o >> 256; o5_X = reg_o; operation : -s*b + a + acc;
"000000100001111000010011000000100000011010110110101110",
--  (2243) addition_subtraction_with_reduction_112
-- reg_a = o6_X; reg_b = 2prime6; reg_acc = reg_o >> 256; o6_X = reg_o; operation : -s*b + a + acc;
"000000100001111000010011000000100000011111011011001110",
--  (2244) addition_subtraction_with_reduction_113
-- reg_a = o7_X; reg_b = 2prime7; reg_acc = reg_o >> 256; o7_X = reg_o; Enable sign a,b; operation : -s*b + a + acc;
"000000100001111000010011000000100001100011111111101110",
--  (2245) addition_subtraction_with_reduction_114
-- reg_a = o0_X; reg_b = 2prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc;
"000000100001111000010001010011010000000100000000001110",
--  (2246) addition_subtraction_with_reduction_115
-- reg_a = o1_X; reg_b = 2prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : s*b + a + acc;
"000000100001111000010001010000100000001000100100101110",
--  (2247) addition_subtraction_with_reduction_116
-- reg_a = o2_X; reg_b = 2prime2; reg_acc = reg_o >> 256; o2_X = reg_o; operation : s*b + a + acc;
"000000100001111000010001010000100000001101001001001110",
--  (2248) addition_subtraction_with_reduction_117
-- reg_a = o3_X; reg_b = 2prime3; reg_acc = reg_o >> 256; o3_X = reg_o; operation : s*b + a + acc;
"000000100001111000010001010000100000010001101101101110",
--  (2249) addition_subtraction_with_reduction_118
-- reg_a = o4_X; reg_b = 2prime4; reg_acc = reg_o >> 256; o4_X = reg_o; operation : s*b + a + acc;
"000000100001111000010001010000100000010110010010001101",
--  (2250) addition_subtraction_with_reduction_119
-- reg_a = o5_X; reg_b = 2prime5; reg_acc = reg_o >> 256; o5_X = reg_o; operation : s*b + a + acc;
"000000100001111000010001010000100000011010110110101110",
--  (2251) addition_subtraction_with_reduction_120
-- reg_a = o6_X; reg_b = 2prime6; reg_acc = reg_o >> 256; o6_X = reg_o; operation : s*b + a + acc;
"000000100001111000010001010000100000011111011011001110",
--  (2252) addition_subtraction_with_reduction_121
-- reg_a = o7_X; reg_b = 2prime7; reg_acc = reg_o >> 256; o7_X = reg_o; Enable sign a,b; operation : s*b + a + acc;
"000000100001111000010001010000100001100011111111101110",
--  (2253) addition_subtraction_with_reduction_122
-- reg_a = o0_X; reg_b = 2prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc;
"000000100001111000010001010011010000000100000000001110",
--  (2254) addition_subtraction_with_reduction_123
-- reg_a = o1_X; reg_b = 2prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : s*b + a + acc;
"000000100001111000010001010000100000001000100100101110",
--  (2255) addition_subtraction_with_reduction_124
-- reg_a = o2_X; reg_b = 2prime2; reg_acc = reg_o >> 256; o2_X = reg_o; operation : s*b + a + acc;
"000000100001111000010001010000100000001101001001001110",
--  (2256) addition_subtraction_with_reduction_125
-- reg_a = o3_X; reg_b = 2prime3; reg_acc = reg_o >> 256; o3_X = reg_o; operation : s*b + a + acc;
"000000100001111000010001010000100000010001101101101110",
--  (2257) addition_subtraction_with_reduction_126
-- reg_a = o4_X; reg_b = 2prime4; reg_acc = reg_o >> 256; o4_X = reg_o; operation : s*b + a + acc;
"000000100001111000010001010000100000010110010010001110",
--  (2258) addition_subtraction_with_reduction_127
-- reg_a = o5_X; reg_b = 2prime5; reg_acc = reg_o >> 256; o5_X = reg_o; operation : s*b + a + acc;
"000000100001111000010001010000100000011010110110101110",
--  (2259) addition_subtraction_with_reduction_128
-- reg_a = o6_X; reg_b = 2prime6; reg_acc = reg_o >> 256; o6_X = reg_o; operation : s*b + a + acc;
"000000100001111000010001010000100000011111011011001110",
--  (2260) addition_subtraction_with_reduction_129
-- reg_a = o7_X; reg_b = 2prime7; reg_acc = reg_o >> 256; o7_X = reg_o; Enable sign a,b; operation : s*b + a + acc;
"000000100001111000010001010000100001100011111111101110",
--  (2261) addition_subtraction_with_reduction_130
-- NOP 4 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : b + a + acc;
"000000000000000100000000010000011110000100000000000010"
);



constant rom_state_machine_fill_nop : romtype(2262 to 4095) := (others => "000000000000000100000000100000011110000100000000000011");
constant rom_state_machine : romtype(0 to 4095) := rom_state_machine_program & rom_state_machine_fill_nop;

signal rom_state_machine_address : std_logic_vector(11 downto 0);
signal rom_state_machine_output : std_logic_vector(53 downto 0);

signal rom_sm_rotation_size : std_logic_vector(1 downto 0);
signal rom_sel_address_a : std_logic;
signal rom_sel_address_b_prime : std_logic_vector(1 downto 0);
signal rom_sm_specific_mac_address_a : std_logic_vector(2 downto 0);
signal rom_sm_specific_mac_address_b : std_logic_vector(2 downto 0);
signal rom_sm_specific_mac_address_o : std_logic_vector(2 downto 0);
signal rom_sm_specific_mac_next_address_o : std_logic_vector(2 downto 0);
signal rom_mac_enable_signed_a : std_logic;
signal rom_mac_enable_signed_b : std_logic;
signal rom_mac_sel_load_reg_a : std_logic_vector(1 downto 0);
signal rom_mac_clear_reg_b : std_logic;
signal rom_mac_clear_reg_acc : std_logic;
signal rom_mac_sel_shift_reg_o : std_logic;
signal rom_mac_enable_update_reg_s : std_logic;
signal rom_mac_sel_reg_s_reg_o_sign : std_logic;
signal rom_mac_reg_s_reg_o_positive : std_logic;
signal rom_sm_sign_a_mode : std_logic;
signal rom_sm_mac_operation_mode : std_logic_vector(1 downto 0);
signal rom_mac_enable_reg_s_mask : std_logic;
signal rom_mac_subtraction_reg_a_b : std_logic;
signal rom_mac_sel_multiply_two_a_b : std_logic;
signal rom_mac_sel_reg_y_output : std_logic;
signal rom_sm_mac_write_enable_output : std_logic;
signal rom_mac_memory_double_mode : std_logic;
signal rom_mac_memory_only_write_mode : std_logic;
signal rom_base_address_generator_o_increment_previous_address : std_logic;

signal rom_last_state : std_logic;
signal rom_current_operand_size : std_logic_vector(2 downto 0);
signal rom_next_operation_same_operand_size : std_logic_vector(4 downto 0);
signal rom_next_operation_different_operand_size : std_logic_vector(6 downto 0);

signal adder_a : unsigned(11 downto 0);
signal adder_b : unsigned(6 downto 0);
signal adder_o : unsigned(11 downto 0);

signal ultimate_instruction : std_logic;

signal internal_sel_output_rom : std_logic;
signal internal_update_rom_address : std_logic;
signal internal_sel_load_new_rom_address : std_logic;
signal internal_sm_rotation_size : std_logic_vector(1 downto 0);
signal internal_sm_circular_shift_enable : std_logic;
signal internal_sel_address_a : std_logic;
signal internal_sel_address_b_prime : std_logic_vector(1 downto 0);
signal internal_sm_specific_mac_address_a : std_logic_vector(2 downto 0);
signal internal_sm_specific_mac_address_b : std_logic_vector(2 downto 0);
signal internal_sm_specific_mac_address_o : std_logic_vector(2 downto 0);
signal internal_sm_specific_mac_next_address_o : std_logic_vector(2 downto 0);
signal internal_mac_enable_signed_a : std_logic;
signal internal_mac_enable_signed_b : std_logic;
signal internal_mac_sel_load_reg_a : std_logic_vector(1 downto 0);
signal internal_mac_clear_reg_b : std_logic;
signal internal_mac_clear_reg_acc : std_logic;
signal internal_mac_sel_shift_reg_o : std_logic;
signal internal_mac_enable_update_reg_s : std_logic;
signal internal_mac_sel_reg_s_reg_o_sign : std_logic;
signal internal_mac_reg_s_reg_o_positive : std_logic;
signal internal_sm_sign_a_mode : std_logic;
signal internal_sm_mac_operation_mode : std_logic_vector(1 downto 0);
signal internal_mac_enable_reg_s_mask : std_logic;
signal internal_mac_subtraction_reg_a_b : std_logic;
signal internal_mac_sel_multiply_two_a_b : std_logic;
signal internal_mac_sel_reg_y_output : std_logic;
signal internal_sm_mac_write_enable_output : std_logic;
signal internal_mac_memory_double_mode : std_logic;
signal internal_mac_memory_only_write_mode : std_logic;
signal internal_base_address_generator_o_increment_previous_address : std_logic;
signal internal_sm_free_flag : std_logic;

-- 0000 multiplication with no reduction
constant first_state_multiplication_direct_operand_size_1 : std_logic_vector(11 downto 0)                                      := std_logic_vector(to_unsigned(0,12));
constant first_state_multiplication_direct_operand_size_2_3_4_5_6_7_8 : std_logic_vector(11 downto 0)                          := std_logic_vector(to_unsigned(2,12));
-- 0001 square with no reduction                                                                                               
constant first_state_square_direct_operand_size_1 : std_logic_vector(11 downto 0)                                              := std_logic_vector(to_unsigned(141,12));
constant first_state_square_direct_operand_size_2_3_4_5_6_7_8 : std_logic_vector(11 downto 0)                                  := std_logic_vector(to_unsigned(143,12));
-- 0010 multiplication with reduction and prime line not equal to 1                                                            
constant first_state_multiplication_with_reduction_operand_size_1 : std_logic_vector(11 downto 0)                              := std_logic_vector(to_unsigned(226,12));
constant first_state_multiplication_with_reduction_operand_size_2_3_4_5_6_7_8 : std_logic_vector(11 downto 0)                  := std_logic_vector(to_unsigned(231,12));
-- 0010 multiplication with reduction and prime line equal to 1                                                     
constant first_state_multiplication_with_reduction_special_prime_1_operand_size_1 : std_logic_vector(11 downto 0)              := std_logic_vector(to_unsigned(510,12));
constant first_state_multiplication_with_reduction_special_prime_1_operand_size_2_3_4_5_6_7_8 : std_logic_vector(11 downto 0)  := std_logic_vector(to_unsigned(513,12));
constant first_state_multiplication_with_reduction_special_prime_2_operand_size_2_3_4_5_6_7_8 : std_logic_vector(11 downto 0)  := std_logic_vector(to_unsigned(765,12));
constant first_state_multiplication_with_reduction_special_prime_3_operand_size_3_4_5_6_7_8 : std_logic_vector(11 downto 0)    := std_logic_vector(to_unsigned(1002,12));
-- 0011 square with reduction and prime line not equal to 1                                                                    
constant first_state_square_with_reduction_operand_size_1 : std_logic_vector(11 downto 0)                                      := std_logic_vector(to_unsigned(1217,12));
constant first_state_square_with_reduction_operand_size_2_3_4_5_6_7_8 : std_logic_vector(11 downto 0)                          := std_logic_vector(to_unsigned(1222,12));
-- 0011 square with reduction and prime line equal to 1                                                                        
constant first_state_square_with_reduction_special_prime_1_operand_size_1 : std_logic_vector(11 downto 0)                      := std_logic_vector(to_unsigned(1445,12));
constant first_state_square_with_reduction_special_prime_1_operand_size_2_3_4_5_6_7_8 : std_logic_vector(11 downto 0)          := std_logic_vector(to_unsigned(1448,12));
constant first_state_square_with_reduction_special_prime_2_operand_size_2_3_4_5_6_7_8 : std_logic_vector(11 downto 0)          := std_logic_vector(to_unsigned(1643,12));
constant first_state_square_with_reduction_special_prime_3_operand_size_3_4_5_6_7_8 : std_logic_vector(11 downto 0)            := std_logic_vector(to_unsigned(1824,12));
-- 0100 addition with no reduction                                                                                             
constant first_state_addition_subtraction_direct_operand_size_1 : std_logic_vector(11 downto 0)                                := std_logic_vector(to_unsigned(1984, 12));
constant first_state_addition_subtraction_direct_operand_size_2_3_4_5_6_7_8 : std_logic_vector(11 downto 0)                    := std_logic_vector(to_unsigned(1986, 12));
-- 0101 iterative modular reduction                                                                                            
constant first_state_iterative_modular_reduction_operand_size_1 : std_logic_vector(11 downto 0)                                := std_logic_vector(to_unsigned(2007, 12));
constant first_state_iterative_modular_reduction_operand_size_2 : std_logic_vector(11 downto 0)                                := std_logic_vector(to_unsigned(2012, 12));
constant first_state_iterative_modular_reduction_operand_size_3 : std_logic_vector(11 downto 0)                                := std_logic_vector(to_unsigned(2020, 12));
constant first_state_iterative_modular_reduction_operand_size_4 : std_logic_vector(11 downto 0)                                := std_logic_vector(to_unsigned(2031, 12));
constant first_state_iterative_modular_reduction_operand_size_5 : std_logic_vector(11 downto 0)                                := std_logic_vector(to_unsigned(2045, 12));
constant first_state_iterative_modular_reduction_operand_size_6 : std_logic_vector(11 downto 0)                                := std_logic_vector(to_unsigned(2062, 12));
constant first_state_iterative_modular_reduction_operand_size_7 : std_logic_vector(11 downto 0)                                := std_logic_vector(to_unsigned(2082, 12));
constant first_state_iterative_modular_reduction_operand_size_8 : std_logic_vector(11 downto 0)                                := std_logic_vector(to_unsigned(2105, 12));
-- 0110 addition with no reduction                                                                                             
constant first_state_addition_subtraction_with_reduction_operand_size_1 : std_logic_vector(11 downto 0)                        := std_logic_vector(to_unsigned(2131, 12));
constant first_state_addition_subtraction_with_reduction_operand_size_2_3_4_5_6_7_8 : std_logic_vector(11 downto 0)            := std_logic_vector(to_unsigned(2136, 12));

type state is (reset, decode_instruction, instruction_execution);

signal actual_state, next_state : state;

signal internal_next_sel_output_rom : std_logic;
signal internal_next_update_rom_address : std_logic;
signal internal_next_sel_load_new_rom_address : std_logic;
signal internal_next_sm_rotation_size : std_logic_vector(1 downto 0);
signal internal_next_sm_circular_shift_enable : std_logic;
signal internal_next_sel_address_a : std_logic;
signal internal_next_sel_address_b_prime : std_logic_vector(1 downto 0);
signal internal_next_sm_specific_mac_address_a : std_logic_vector(2 downto 0);
signal internal_next_sm_specific_mac_address_b : std_logic_vector(2 downto 0);
signal internal_next_sm_specific_mac_address_o : std_logic_vector(2 downto 0);
signal internal_next_sm_specific_mac_next_address_o : std_logic_vector(2 downto 0);
signal internal_next_mac_enable_signed_a : std_logic;
signal internal_next_mac_enable_signed_b : std_logic;
signal internal_next_mac_sel_load_reg_a : std_logic_vector(1 downto 0);
signal internal_next_mac_clear_reg_b : std_logic;
signal internal_next_mac_clear_reg_acc : std_logic;
signal internal_next_mac_sel_shift_reg_o : std_logic;
signal internal_next_mac_enable_update_reg_s : std_logic;
signal internal_next_mac_sel_reg_s_reg_o_sign : std_logic;
signal internal_next_mac_reg_s_reg_o_positive : std_logic;
signal internal_next_sm_sign_a_mode : std_logic;
signal internal_next_sm_mac_operation_mode : std_logic_vector(1 downto 0);
signal internal_next_mac_enable_reg_s_mask : std_logic;
signal internal_next_mac_subtraction_reg_a_b : std_logic;
signal internal_next_mac_sel_multiply_two_a_b : std_logic;
signal internal_next_mac_sel_reg_y_output : std_logic;
signal internal_next_sm_mac_write_enable_output : std_logic;
signal internal_next_mac_memory_double_mode : std_logic;
signal internal_next_mac_memory_only_write_mode : std_logic;
signal internal_next_base_address_generator_o_increment_previous_address : std_logic;
signal internal_next_sm_free_flag : std_logic;

begin

registers_state : process(clk, rstn)
begin
    if(rstn = '0') then
        actual_state <= reset;
    elsif(rising_edge(clk)) then
        actual_state <= next_state;
    end if;
end process;

registers_state_output : process(clk)
begin
    if(rising_edge(clk)) then
        if(rstn = '0') then
            internal_sel_output_rom <= '0';
            internal_update_rom_address <= '1';
            internal_sel_load_new_rom_address <= '1';
            internal_sm_rotation_size <= "11";
            internal_sm_circular_shift_enable <= '0';
            internal_sel_address_a <= '0';
            internal_sel_address_b_prime <= "00";
            internal_sm_specific_mac_address_a <= "000";
            internal_sm_specific_mac_address_b <= "000";
            internal_sm_specific_mac_address_o <= "000";
            internal_sm_specific_mac_next_address_o <= "001";
            internal_mac_enable_signed_a <= '0';
            internal_mac_enable_signed_b <= '0';
            internal_mac_sel_load_reg_a <= "00";
            internal_mac_clear_reg_b <= '0';
            internal_mac_clear_reg_acc <= '0';
            internal_mac_sel_shift_reg_o <= '0';
            internal_mac_enable_update_reg_s <= '0';
            internal_mac_sel_reg_s_reg_o_sign <= '0';
            internal_mac_reg_s_reg_o_positive <= '0';
            internal_sm_sign_a_mode <= '0';
            internal_sm_mac_operation_mode <= "00";
            internal_mac_enable_reg_s_mask <= '0';
            internal_mac_subtraction_reg_a_b <= '0';
            internal_mac_sel_multiply_two_a_b <= '0';
            internal_mac_sel_reg_y_output <= '0';
            internal_sm_mac_write_enable_output <= '0';
            internal_mac_memory_double_mode <= '0';
            internal_mac_memory_only_write_mode <= '0';
            internal_base_address_generator_o_increment_previous_address <= '0';
            internal_sm_free_flag <= '0';
        else
            internal_sel_output_rom <= internal_next_sel_output_rom;
            internal_update_rom_address <= internal_next_update_rom_address;
            internal_sel_load_new_rom_address <= internal_next_sel_load_new_rom_address;
            internal_sm_rotation_size <= internal_next_sm_rotation_size;
            internal_sm_circular_shift_enable <= internal_next_sm_circular_shift_enable;
            internal_sel_address_a <= internal_next_sel_address_a;
            internal_sel_address_b_prime <= internal_next_sel_address_b_prime;
            internal_sm_specific_mac_address_a <= internal_next_sm_specific_mac_address_a;
            internal_sm_specific_mac_address_b <= internal_next_sm_specific_mac_address_b;
            internal_sm_specific_mac_address_o <= internal_next_sm_specific_mac_address_o;
            internal_sm_specific_mac_next_address_o <= internal_next_sm_specific_mac_next_address_o;
            internal_mac_enable_signed_a <= internal_next_mac_enable_signed_a;
            internal_mac_enable_signed_b <= internal_next_mac_enable_signed_b;
            internal_mac_sel_load_reg_a <= internal_next_mac_sel_load_reg_a;
            internal_mac_clear_reg_b <= internal_next_mac_clear_reg_b;
            internal_mac_clear_reg_acc <= internal_next_mac_clear_reg_acc;
            internal_mac_sel_shift_reg_o <= internal_next_mac_sel_shift_reg_o;
            internal_mac_enable_update_reg_s <= internal_next_mac_enable_update_reg_s;
            internal_mac_sel_reg_s_reg_o_sign <= internal_next_mac_sel_reg_s_reg_o_sign;
            internal_mac_reg_s_reg_o_positive <= internal_next_mac_reg_s_reg_o_positive;
            internal_sm_sign_a_mode <= internal_next_sm_sign_a_mode;
            internal_sm_mac_operation_mode <= internal_next_sm_mac_operation_mode;
            internal_mac_enable_reg_s_mask <= internal_next_mac_enable_reg_s_mask;
            internal_mac_subtraction_reg_a_b <= internal_next_mac_subtraction_reg_a_b;
            internal_mac_sel_multiply_two_a_b <= internal_next_mac_sel_multiply_two_a_b;
            internal_mac_sel_reg_y_output <= internal_next_mac_sel_reg_y_output;
            internal_sm_mac_write_enable_output <= internal_next_sm_mac_write_enable_output;
            internal_mac_memory_double_mode <= internal_next_mac_memory_double_mode;
            internal_mac_memory_only_write_mode <= internal_next_mac_memory_only_write_mode;
            internal_base_address_generator_o_increment_previous_address <= internal_next_base_address_generator_o_increment_previous_address;
            internal_sm_free_flag <= internal_next_sm_free_flag;
        end if;
    end if;
end process;

update_output : process(actual_state, instruction_values_valid, instruction_type)
begin
    case (actual_state) is
        when reset =>
            internal_next_sel_output_rom <= '0';
            internal_next_update_rom_address <= '1';
            internal_next_sel_load_new_rom_address <= '1';
            internal_next_sm_rotation_size <= "11";
            internal_next_sm_circular_shift_enable <= '0';
            internal_next_sel_address_a <= '0';
            internal_next_sel_address_b_prime <= "00";
            internal_next_sm_specific_mac_address_a <= "000";
            internal_next_sm_specific_mac_address_b <= "000";
            internal_next_sm_specific_mac_address_o <= "000";
            internal_next_sm_specific_mac_next_address_o <= "001";
            internal_next_mac_enable_signed_a <= '0';
            internal_next_mac_enable_signed_b <= '0';
            internal_next_mac_sel_load_reg_a <= "11";
            internal_next_mac_clear_reg_b <= '1';
            internal_next_mac_clear_reg_acc <= '1';
            internal_next_mac_sel_shift_reg_o <= '0';
            internal_next_mac_enable_update_reg_s <= '0';
            internal_next_mac_sel_reg_s_reg_o_sign <= '0';
            internal_next_mac_reg_s_reg_o_positive <= '0';
            internal_next_sm_sign_a_mode <= '0';
            internal_next_sm_mac_operation_mode <= "10";
            internal_next_mac_enable_reg_s_mask <= '0';
            internal_next_mac_subtraction_reg_a_b <= '0';
            internal_next_mac_sel_multiply_two_a_b <= '0';
            internal_next_mac_sel_reg_y_output <= '0';
            internal_next_sm_mac_write_enable_output <= '0';
            internal_next_mac_memory_double_mode <= '0';
            internal_next_mac_memory_only_write_mode <= '0';
            internal_next_base_address_generator_o_increment_previous_address <= '0';
            internal_next_sm_free_flag <= '1';
        when decode_instruction =>
            internal_next_sel_output_rom <= '0';
            internal_next_update_rom_address <= '1';
            internal_next_sel_load_new_rom_address <= '1';
            internal_next_sm_free_flag <= '1';
            internal_next_sm_rotation_size <= "11";
            internal_next_sm_circular_shift_enable <= '0';
            internal_next_sel_address_a <= '0';
            internal_next_sel_address_b_prime <= "00";
            internal_next_sm_specific_mac_address_a <= "000";
            internal_next_sm_specific_mac_address_b <= "000";
            internal_next_sm_specific_mac_address_o <= "000";
            internal_next_sm_specific_mac_next_address_o <= "001";
            internal_next_mac_enable_signed_a <= '0';
            internal_next_mac_enable_signed_b <= '0';
            internal_next_mac_sel_load_reg_a <= "11";
            internal_next_mac_clear_reg_b <= '1';
            internal_next_mac_clear_reg_acc <= '1';
            internal_next_mac_sel_shift_reg_o <= '0';
            internal_next_mac_enable_update_reg_s <= '0';
            internal_next_mac_sel_reg_s_reg_o_sign <= '0';
            internal_next_mac_reg_s_reg_o_positive <= '0';
            internal_next_sm_sign_a_mode <= '0';
            internal_next_sm_mac_operation_mode <= "10";
            internal_next_mac_enable_reg_s_mask <= '0';
            internal_next_mac_subtraction_reg_a_b <= '0';
            internal_next_mac_sel_multiply_two_a_b <= '0';
            internal_next_mac_sel_reg_y_output <= '0';
            internal_next_sm_mac_write_enable_output <= '0';
            internal_next_mac_memory_double_mode <= '0';
            internal_next_mac_memory_only_write_mode <= '0';
            internal_next_base_address_generator_o_increment_previous_address <= '0';
            if(instruction_values_valid = '1') then
                internal_next_sm_free_flag <= '0';
                internal_next_sel_output_rom <= '1';
                internal_next_update_rom_address <= '1';
                internal_next_sel_load_new_rom_address <= '0';
                internal_next_sm_free_flag <= '0';
                internal_next_sm_circular_shift_enable <= '1';
                if(instruction_type = "0000") then
                    internal_next_sm_rotation_size <= "11";
                elsif(instruction_type = "0001") then
                    internal_next_sm_rotation_size <= "11";
                elsif(instruction_type = "0010") then
                    internal_next_sm_rotation_size <= "11";
                elsif(instruction_type = "0011") then
                    internal_next_sm_rotation_size <= "11";
                elsif(instruction_type = "0100") then
                    internal_next_sm_rotation_size <= "10";
                elsif(instruction_type = "0101") then
                    internal_next_sm_rotation_size <= "10";
                elsif(instruction_type = "0110") then
                    internal_next_sm_rotation_size <= "10";
                end if;
            end if;
        when instruction_execution =>
            internal_next_sel_output_rom <= '1';
            internal_next_update_rom_address <= '1';
            internal_next_sel_load_new_rom_address <= '0';
            internal_next_sm_free_flag <= '0';
            internal_next_sm_rotation_size <= "11";
            internal_next_sm_circular_shift_enable <= '1';
            internal_next_sel_address_a <= '0';
            internal_next_sel_address_b_prime <= "00";
            internal_next_sm_specific_mac_address_a <= "000";
            internal_next_sm_specific_mac_address_b <= "000";
            internal_next_sm_specific_mac_address_o <= "000";
            internal_next_sm_specific_mac_next_address_o <= "001";
            internal_next_mac_enable_signed_a <= '0';
            internal_next_mac_enable_signed_b <= '0';
            internal_next_mac_sel_load_reg_a <= "11";
            internal_next_mac_clear_reg_b <= '1';
            internal_next_mac_clear_reg_acc <= '1';
            internal_next_mac_sel_shift_reg_o <= '0';
            internal_next_mac_enable_update_reg_s <= '0';
            internal_next_mac_sel_reg_s_reg_o_sign <= '0';
            internal_next_mac_reg_s_reg_o_positive <= '0';
            internal_next_sm_sign_a_mode <= '0';
            internal_next_sm_mac_operation_mode <= "10";
            internal_next_mac_enable_reg_s_mask <= '0';
            internal_next_mac_subtraction_reg_a_b <= '0';
            internal_next_mac_sel_multiply_two_a_b <= '0';
            internal_next_mac_sel_reg_y_output <= '0';
            internal_next_sm_mac_write_enable_output <= '0';
            internal_next_mac_memory_double_mode <= '0';
            internal_next_mac_memory_only_write_mode <= '0';
            internal_next_base_address_generator_o_increment_previous_address <= '0';
    end case;
end process;

update_state : process(actual_state, instruction_type, operands_size, instruction_values_valid, penultimate_operation, rom_last_state)
begin
case (actual_state) is
        when reset =>
            next_state <= decode_instruction;
        when decode_instruction =>
            next_state <= decode_instruction;
            if(instruction_values_valid = '1') then
                next_state <= instruction_execution;
            end if;
        when instruction_execution =>
            next_state <= instruction_execution;
            if((penultimate_operation = '1') and (rom_last_state = '1')) then
                next_state <= decode_instruction;
            end if;
end case;
end process;

process(clk)
begin
    if(rising_edge(clk)) then
        if(rstn = '0') then
            ultimate_instruction <= '0';
        else
            ultimate_instruction <= penultimate_operation;
        end if;
    end if;
end process;

adder_a <= unsigned(rom_state_machine_address);
adder_b <= resize(unsigned(rom_next_operation_same_operand_size), adder_b'length) when (rom_current_operand_size = operands_size) else unsigned(rom_next_operation_different_operand_size);

adder_o <= adder_a + resize(adder_b, adder_o'length);

process(clk)
begin
    if (rising_edge(clk)) then
        if(internal_update_rom_address = '1') then
            if(internal_sel_load_new_rom_address = '1') then
                if(instruction_values_valid = '1') then
                    if(instruction_type = "0000") then
                        if(operands_size = "000") then
                            rom_state_machine_address <= first_state_multiplication_direct_operand_size_1;
                        else
                            rom_state_machine_address <= first_state_multiplication_direct_operand_size_2_3_4_5_6_7_8;
                        end if;
                    elsif(instruction_type = "0001") then
                        if(operands_size = "000") then
                            rom_state_machine_address <= first_state_square_direct_operand_size_1;
                        else
                            rom_state_machine_address <= first_state_square_direct_operand_size_2_3_4_5_6_7_8;
                        end if;
                    elsif(instruction_type = "0010") then
                        case (prime_line_equal_one) is
                            when "00" =>
                                if(operands_size = "000") then
                                    rom_state_machine_address <= first_state_multiplication_with_reduction_operand_size_1;
                                else
                                    rom_state_machine_address <= first_state_multiplication_with_reduction_operand_size_2_3_4_5_6_7_8;
                                end if;
                            when "01" =>
                                if(operands_size = "000") then
                                    rom_state_machine_address <= first_state_multiplication_with_reduction_special_prime_1_operand_size_1;
                                else
                                    rom_state_machine_address <= first_state_multiplication_with_reduction_special_prime_1_operand_size_2_3_4_5_6_7_8;
                                end if;
                            when "10" =>
                                rom_state_machine_address <= first_state_multiplication_with_reduction_special_prime_2_operand_size_2_3_4_5_6_7_8;
                            when "11" =>
                                rom_state_machine_address <= first_state_multiplication_with_reduction_special_prime_3_operand_size_3_4_5_6_7_8;
                            when others =>
                                rom_state_machine_address <= std_logic_vector(to_unsigned(0, rom_state_machine_address'length));
                        end case;
                    elsif(instruction_type = "0011") then
                        case (prime_line_equal_one) is
                            when "00" =>
                                if(operands_size = "000") then
                                    rom_state_machine_address <= first_state_square_with_reduction_operand_size_1;
                                else
                                    rom_state_machine_address <= first_state_square_with_reduction_operand_size_2_3_4_5_6_7_8;
                                end if;
                            when "01" =>
                                if(operands_size = "000") then
                                    rom_state_machine_address <= first_state_square_with_reduction_special_prime_1_operand_size_1;
                                else
                                    rom_state_machine_address <= first_state_square_with_reduction_special_prime_1_operand_size_2_3_4_5_6_7_8;
                                end if;
                            when "10" =>
                                rom_state_machine_address <= first_state_square_with_reduction_special_prime_2_operand_size_2_3_4_5_6_7_8;
                            when "11" =>
                                rom_state_machine_address <= first_state_square_with_reduction_special_prime_3_operand_size_3_4_5_6_7_8;
                            when others =>
                                rom_state_machine_address <= std_logic_vector(to_unsigned(0, rom_state_machine_address'length));
                        end case;
                    elsif(instruction_type = "0100") then
                        if(operands_size = "000") then
                            rom_state_machine_address <= first_state_addition_subtraction_direct_operand_size_1;
                        else
                            rom_state_machine_address <= first_state_addition_subtraction_direct_operand_size_2_3_4_5_6_7_8;
                        end if;
                    elsif(instruction_type = "0101") then
                        if(operands_size = "000") then
                            rom_state_machine_address <= first_state_iterative_modular_reduction_operand_size_1;
                        elsif(operands_size = "001") then
                            rom_state_machine_address <= first_state_iterative_modular_reduction_operand_size_2;
                        elsif(operands_size = "010") then
                            rom_state_machine_address <= first_state_iterative_modular_reduction_operand_size_3;
                        elsif(operands_size = "011") then
                            rom_state_machine_address <= first_state_iterative_modular_reduction_operand_size_4;
                        elsif(operands_size = "100") then
                            rom_state_machine_address <= first_state_iterative_modular_reduction_operand_size_5;
                        elsif(operands_size = "101") then
                            rom_state_machine_address <= first_state_iterative_modular_reduction_operand_size_6;
                        elsif(operands_size = "110") then
                            rom_state_machine_address <= first_state_iterative_modular_reduction_operand_size_7;
                        else
                            rom_state_machine_address <= first_state_iterative_modular_reduction_operand_size_8;
                        end if;
                    elsif(instruction_type = "0110") then
                        if(operands_size = "000") then
                            rom_state_machine_address <= first_state_addition_subtraction_with_reduction_operand_size_1;
                        else
                            rom_state_machine_address <= first_state_addition_subtraction_with_reduction_operand_size_2_3_4_5_6_7_8;
                        end if;
                    end if;
                end if;
            elsif(ultimate_instruction = '1') then
                rom_state_machine_address <= std_logic_vector(adder_o);
            end if;
        end if;
    end if;
end process;

rom_state_machine_output <= rom_state_machine(to_integer(to_01(unsigned(rom_state_machine_address))));

rom_sm_rotation_size <= rom_state_machine_output(1 downto 0);
rom_sel_address_a <= rom_state_machine_output(2);
rom_sel_address_b_prime <= rom_state_machine_output(4 downto 3);
rom_sm_specific_mac_address_a <= rom_state_machine_output(7 downto 5);
rom_sm_specific_mac_address_b <= rom_state_machine_output(10 downto 8);
rom_sm_specific_mac_address_o <= rom_state_machine_output(13 downto 11);
rom_sm_specific_mac_next_address_o <= rom_state_machine_output(16 downto 14);
rom_mac_enable_signed_a <= rom_state_machine_output(17);
rom_mac_enable_signed_b <= rom_state_machine_output(18);
rom_mac_sel_load_reg_a <= rom_state_machine_output(20 downto 19);
rom_mac_clear_reg_b <= rom_state_machine_output(21);
rom_mac_clear_reg_acc <= rom_state_machine_output(22);
rom_mac_sel_shift_reg_o <= rom_state_machine_output(23);
rom_mac_enable_update_reg_s <= rom_state_machine_output(24);
rom_mac_sel_reg_s_reg_o_sign <= rom_state_machine_output(25);
rom_mac_reg_s_reg_o_positive <= rom_state_machine_output(26);
rom_sm_sign_a_mode <= rom_state_machine_output(27);
rom_sm_mac_operation_mode <= rom_state_machine_output(29 downto 28);
rom_mac_enable_reg_s_mask <= rom_state_machine_output(30);
rom_mac_subtraction_reg_a_b <= rom_state_machine_output(31);
rom_mac_sel_multiply_two_a_b <= rom_state_machine_output(32);
rom_mac_sel_reg_y_output <= rom_state_machine_output(33);
rom_sm_mac_write_enable_output <= rom_state_machine_output(34);
rom_mac_memory_double_mode <= rom_state_machine_output(35);
rom_mac_memory_only_write_mode <= rom_state_machine_output(36);
rom_base_address_generator_o_increment_previous_address <= rom_state_machine_output(37);

rom_last_state <= rom_state_machine_output(38);
rom_current_operand_size <= rom_state_machine_output(41 downto 39);
rom_next_operation_same_operand_size <= rom_state_machine_output(46 downto 42);
rom_next_operation_different_operand_size <= rom_state_machine_output(53 downto 47);

sm_rotation_size <= rom_sm_rotation_size when internal_sel_output_rom = '1' else internal_sm_rotation_size;
sm_circular_shift_enable <= internal_sm_circular_shift_enable;
sel_address_a <= rom_sel_address_a when internal_sel_output_rom = '1' else internal_sel_address_a;
sel_address_b_prime <= rom_sel_address_b_prime when internal_sel_output_rom = '1' else internal_sel_address_b_prime;
sm_specific_mac_address_a <= rom_sm_specific_mac_address_a when internal_sel_output_rom = '1' else internal_sm_specific_mac_address_a;
sm_specific_mac_address_b <= rom_sm_specific_mac_address_b when internal_sel_output_rom = '1' else internal_sm_specific_mac_address_b;
sm_specific_mac_address_o <= rom_sm_specific_mac_address_o when internal_sel_output_rom = '1' else internal_sm_specific_mac_address_o;
sm_specific_mac_next_address_o <= rom_sm_specific_mac_next_address_o when internal_sel_output_rom = '1' else internal_sm_specific_mac_next_address_o;
mac_enable_signed_a <= rom_mac_enable_signed_a when internal_sel_output_rom = '1' else internal_mac_enable_signed_a;
mac_enable_signed_b <= rom_mac_enable_signed_b when internal_sel_output_rom = '1' else internal_mac_enable_signed_b;
mac_sel_load_reg_a <= rom_mac_sel_load_reg_a when internal_sel_output_rom = '1' else internal_mac_sel_load_reg_a;
mac_clear_reg_b <= rom_mac_clear_reg_b when internal_sel_output_rom = '1' else internal_mac_clear_reg_b;
mac_clear_reg_acc <= rom_mac_clear_reg_acc when internal_sel_output_rom = '1' else internal_mac_clear_reg_acc;
mac_sel_shift_reg_o <= rom_mac_sel_shift_reg_o when internal_sel_output_rom = '1' else internal_mac_sel_shift_reg_o;
mac_enable_update_reg_s <= rom_mac_enable_update_reg_s when internal_sel_output_rom = '1' else internal_mac_enable_update_reg_s;
mac_sel_reg_s_reg_o_sign <= rom_mac_sel_reg_s_reg_o_sign when internal_sel_output_rom = '1' else internal_mac_sel_reg_s_reg_o_sign;
mac_reg_s_reg_o_positive <= rom_mac_reg_s_reg_o_positive when internal_sel_output_rom = '1' else internal_mac_reg_s_reg_o_positive;
sm_sign_a_mode <= rom_sm_sign_a_mode when internal_sel_output_rom = '1' else internal_sm_sign_a_mode;
sm_mac_operation_mode <= rom_sm_mac_operation_mode when internal_sel_output_rom = '1' else internal_sm_mac_operation_mode;
mac_enable_reg_s_mask <= rom_mac_enable_reg_s_mask when internal_sel_output_rom = '1' else internal_mac_enable_reg_s_mask;
mac_subtraction_reg_a_b <= rom_mac_subtraction_reg_a_b when internal_sel_output_rom = '1' else internal_mac_subtraction_reg_a_b;
mac_sel_multiply_two_a_b <= rom_mac_sel_multiply_two_a_b when internal_sel_output_rom = '1' else internal_mac_sel_multiply_two_a_b;
mac_sel_reg_y_output <= rom_mac_sel_reg_y_output when internal_sel_output_rom = '1' else internal_mac_sel_reg_y_output;
sm_mac_write_enable_output <= rom_sm_mac_write_enable_output when internal_sel_output_rom = '1' else internal_sm_mac_write_enable_output;
mac_memory_double_mode <= rom_mac_memory_double_mode when internal_sel_output_rom = '1' else internal_mac_memory_double_mode;
mac_memory_only_write_mode <= rom_mac_memory_only_write_mode when internal_sel_output_rom = '1' else internal_mac_memory_only_write_mode;
base_address_generator_o_increment_previous_address <= rom_base_address_generator_o_increment_previous_address when internal_sel_output_rom = '1' else internal_base_address_generator_o_increment_previous_address;
sm_free_flag <= internal_sm_free_flag;

end compact_memory_based_v2;







































architecture compact_memory_based_v3 of carmela_state_machine_v128 is

type romtype is array(integer range <>) of std_logic_vector(53 downto 0);

constant rom_state_machine_program : romtype(0 to 2261) := (
--  (0) multiplication_direct_0
-- -- In case of size 1
-- reg_a = a0_X; reg_b = b0_X; reg_acc = 0; o0_X = reg_o; o1_X = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001000001110000100000010001100100000000000011",
--  (1) multiplication_direct_1
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (2) multiplication_direct_2
-- -- Other cases
-- reg_a = a0_X; reg_b = b0_X; reg_acc = 0; o0_X = reg_o; operation : a*b + acc; o0_X = reg_o;
"000010100001001000010000100000010000000100000000000011",
--  (3) multiplication_direct_3
-- -- In case of size 2
-- reg_a = a1_X; reg_b = b0_X; reg_acc = reg_o >> 256; Enable sign a; operation : a*b + acc;
"000000100001001000000000100000100000101000100000100011",
--  (4) multiplication_direct_4
-- reg_a = a0_X; reg_b = b1_X; reg_acc = reg_o; o1_X = reg_o; Enable sign b; operation : a*b + acc;
"000000100001001000010000100000000001001000100100000011",
--  (5) multiplication_direct_5
-- reg_a = a1_X; reg_b = b1_X; reg_acc = reg_o >> 256; o2_X = reg_o; o3_X = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001001001110000100000100000001101000100100011",
--  (6) multiplication_direct_6
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (7) multiplication_direct_7
-- -- Other cases
-- reg_a = a1_X; reg_b = b0_X; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001010000000000100000100000001000100000100011",
--  (8) multiplication_direct_8
-- reg_a = a0_X; reg_b = b1_X; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
"000000100001010000010000100000000000001000100100000011",
--  (9) multiplication_direct_9
-- reg_a = a1_X; reg_b = b1_X; reg_acc = reg_o >> 256; operation : a*b + acc;
"000011100001010000000000100000100000001101000100100011",
--  (10) multiplication_direct_10
-- -- In case of size 3
-- reg_a = a0_X; reg_b = b2_X; reg_acc = reg_o; Enable sign b; operation : a*b + acc;
"000000100001010000000000100000000001001101001000000011",
--  (11) multiplication_direct_11
-- reg_a = a2_X; reg_b = b0_X; reg_acc = reg_o; Enable sign a; o2_X = reg_o; operation : a*b + acc;
"000000100001010000010000100000000000101101000001000011",
--  (12) multiplication_direct_12
-- reg_a = a2_X; reg_b = b1_X; reg_acc = reg_o >> 256; Enable sign a; operation : a*b + acc;
"000000100001010000000000100000100000110001100101000011",
--  (13) multiplication_direct_13
-- reg_a = a1_X; reg_b = b2_X; reg_acc = reg_o; o3_X = reg_o; Enable sign b; operation : a*b + acc;
"000000100001010000010000100000000001010001101000100011",
--  (14) multiplication_direct_14
-- reg_a = a2_X; reg_b = b2_X; reg_acc = reg_o >> 256; o4_X = reg_o; o5_X = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001010001110000100000100001110110001001000011",
--  (15) multiplication_direct_15
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (16) multiplication_direct_16
-- -- Other cases
-- reg_a = a0_0; reg_b = b2_0; reg_acc = reg_o; operation : a*b + acc;
"000000100001011000000000100000000000001101001000000011",
--  (17) multiplication_direct_17
-- reg_a = a2_X; reg_b = b0_X; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
"000000100001011000010000100000000000001101000001000011",
--  (18) multiplication_direct_18
-- reg_a = a2_X; reg_b = b1_X; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001011000000000100000100000010001100101000011",
--  (19) multiplication_direct_19
-- reg_a = a1_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000101000001011000000000100000000000010001101000100011",
--  (20) multiplication_direct_20
-- -- In case of size 4
-- reg_a = a3_X; reg_b = b0_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001011000000000100000000000110001100001100011",
--  (21) multiplication_direct_21
-- reg_a = a0_X; reg_b = b3_X; reg_acc = reg_o; o3_X = reg_o; Enable sign b; operation : a*b + acc;
"000000100001011000010000100000000001010001101100000011",
--  (22) multiplication_direct_22
-- reg_a = a2_X; reg_b = b2_X; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001011000000000100000100000010110001001000011",
--  (23) multiplication_direct_23
-- reg_a = a3_X; reg_b = b1_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001011000000000100000000000110110000101100011",
--  (24) multiplication_direct_24
-- reg_a = a1_X; reg_b = b3_X; reg_acc = reg_o; o4_X = reg_o; Enable sign b; operation : a*b + acc;
"000000100001011000010000100000000001010110001100100011",
--  (25) multiplication_direct_25
-- reg_a = a3_X; reg_b = b2_X; reg_acc = reg_o >> 256; Enable sign a; operation : a*b + acc;
"000000100001011000000000100000100000111010101001100011",
--  (26) multiplication_direct_26
-- reg_a = a2_X; reg_b = b3_X; reg_acc = reg_o; o5_X = reg_o; Enable sign b; operation : a*b + acc;
"000000100001011000010000100000000001011010101101000011",
--  (27) multiplication_direct_27
-- reg_a = a3_X; reg_b = b3_X; reg_acc = reg_o >> 256; o6_X = reg_o; o7_X = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001011001110000100000100001111111001101100011",
--  (28) multiplication_direct_28
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (29) multiplication_direct_29
-- -- Other cases
-- reg_a = a3_X; reg_b = b0_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000010001100001100011",
--  (30) multiplication_direct_30
-- reg_a = a0_X; reg_b = b3_X; reg_acc = reg_o; o3_0 = reg_o; operation : a*b + acc;
"000000100001100000010000100000000000010001101100000011",
--  (31) multiplication_direct_31
-- reg_a = a2_X; reg_b = b2_X; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001100000000000100000100000010110001001000011",
--  (32) multiplication_direct_32
-- reg_a = a3_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000010110000101100011",
--  (33) multiplication_direct_33
-- reg_a = a1_X; reg_b = b3_X; reg_acc = reg_o; o4_0 = reg_o; operation : a*b + acc;
"000111000001100000010000100000000000010110001100100011",
--  (34) multiplication_direct_34
-- -- In case of size 5
-- reg_a = a4_X; reg_b = b0_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001100000000000100000000000110110000010000011",
--  (35) multiplication_direct_35
-- reg_a = a0_X; reg_b = b4_X; reg_acc = reg_o; o4_0 = reg_o; Enable sign b; operation : a*b + acc;
"000000100001100000010000100000000001010110010000000011",
--  (36) multiplication_direct_36
-- reg_a = a3_X; reg_b = b2_X; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001100000000000100000100000011010101001100011",
--  (37) multiplication_direct_37
-- reg_a = a2_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000011010101101000011",
--  (38) multiplication_direct_38
-- reg_a = a4_X; reg_b = b1_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001100000000000100000000000111010100110000011",
--  (39) multiplication_direct_39
-- reg_a = a1_X; reg_b = b4_X; reg_acc = reg_o; o5_X = reg_o; Enable sign b; operation : a*b + acc;
"000000100001100000010000100000000001011010110000100011",
--  (40) multiplication_direct_40
-- reg_a = a3_X; reg_b = b3_X; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001100000000000100000100000011111001101100011",
--  (41) multiplication_direct_41
-- reg_a = a4_X; reg_b = b2_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001100000000000100000000000111111001010000011",
--  (42) multiplication_direct_42
-- reg_a = a2_X; reg_b = b4_X; reg_acc = reg_o; o6_X = reg_o; Enable sign b; operation : a*b + acc;
"000000100001100000010000100000000001011111010001000011",
--  (43) multiplication_direct_43
-- reg_a = a4_X; reg_b = b3_X; reg_acc = reg_o >> 256; Enable sign a; operation : a*b + acc;
"000000100001100000000000100000100000100011101110000011",
--  (44) multiplication_direct_44
-- reg_a = a3_X; reg_b = b4_X; reg_acc = reg_o; o7_X = reg_o; Enable sign b; operation : a*b + acc; Increment base address o;
"000000100001100010010000100000000001000011110001100011",
--  (45) multiplication_direct_45
-- reg_a = a4_X; reg_b = b4_X; reg_acc = reg_o >> 256; o8_X = reg_o; o9_X = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001100001110000100000100001100100010010000011",
--  (46) multiplication_direct_46
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (47) multiplication_direct_47
-- -- Other cases
-- reg_a = a4_X; reg_b = b0_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000010110000010000011",
--  (48) multiplication_direct_48
-- reg_a = a0_X; reg_b = b4_X; reg_acc = reg_o; o4_X = reg_o; operation : a*b + acc;
"000000100001101000010000100000000000010110010000000011",
--  (49) multiplication_direct_49
-- reg_a = a3_X; reg_b = b2_X; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001101000000000100000100000011010101001100011",
--  (50) multiplication_direct_50
-- reg_a = a2_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000011010101101000011",
--  (51) multiplication_direct_51
-- reg_a = a4_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000011010100110000011",
--  (52) multiplication_direct_52
-- reg_a = a1_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"001001100001101000000000100000000000011010110000100011",
--  (53) multiplication_direct_53
-- -- In case of size 6
-- reg_a = a5_X; reg_b = b0_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001101000000000100000000000111010100010100011",
--  (54) multiplication_direct_54
-- reg_a = a0_X; reg_b = b5_X; reg_acc = reg_o; o5_0 = reg_o; Enable sign b; operation : a*b + acc;
"000000100001101000010000100000000001011010110100000011",
--  (55) multiplication_direct_55
-- reg_a = a3_X; reg_b = b3_X; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001101000000000100000100000011111001101100011",
--  (56) multiplication_direct_56
-- reg_a = a2_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000011111010001000011",
--  (57) multiplication_direct_57
-- reg_a = a4_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000011111001010000011",
--  (58) multiplication_direct_58
-- reg_a = a5_X; reg_b = b1_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001101000000000100000000000111111000110100011",
--  (59) multiplication_direct_59
-- reg_a = a1_X; reg_b = b5_X; reg_acc = reg_o; o6_0 = reg_o; Enable sign b; operation : a*b + acc;
"000000100001101000010000100000000001011111010100100011",
--  (60) multiplication_direct_60
-- reg_a = a4_X; reg_b = b3_X; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001101000000000100000100000000011101110000011",
--  (61) multiplication_direct_61
-- reg_a = a3_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000011110001100011",
--  (62) multiplication_direct_62
-- reg_a = a5_X; reg_b = b2_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001101000000000100000000000100011101010100011",
--  (63) multiplication_direct_63
-- reg_a = a2_X; reg_b = b5_X; reg_acc = reg_o; o7_0 = reg_o; Enable sign b; operation : a*b + acc; Increment base address o;
"000000100001101010010000100000000001000011110101000011",
--  (64) multiplication_direct_64
-- reg_a = a4_X; reg_b = b4_X; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001101000000000100000100000000100010010000011",
--  (65) multiplication_direct_65
-- reg_a = a5_X; reg_b = b3_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001101000000000100000000000100100001110100011",
--  (66) multiplication_direct_66
-- reg_a = a3_X; reg_b = b5_X; reg_acc = reg_o; o8_0 = reg_o; Enable sign b; operation : a*b + acc;
"000000100001101000010000100000000001000100010101100011",
--  (67) multiplication_direct_67
-- reg_a = a5_X; reg_b = b4_X; reg_acc = reg_o >> 256; Enable sign a; operation : a*b + acc;
"000000100001101000000000100000100000101000110010100011",
--  (68) multiplication_direct_68
-- reg_a = a4_X; reg_b = b5_X; reg_acc = reg_o; o9_0 = reg_o; Enable sign b; operation : a*b + acc;
"000000100001101000010000100000000001001000110110000011",
--  (69) multiplication_direct_69
-- reg_a = a5_X; reg_b = b5_X; reg_acc = reg_o >> 256; o10_X = reg_o; o11_X = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001101001110000100000100001101101010110100011",
--  (70) multiplication_direct_70
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (71) multiplication_direct_71
-- -- Other cases
-- reg_a = a5_X; reg_b = b0_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000011010100010100011",
--  (72) multiplication_direct_72
-- reg_a = a0_X; reg_b = b5_X; reg_acc = reg_o; o5_0 = reg_o; operation : a*b + acc;
"000000100001110000010000100000000000011010110100000011",
--  (73) multiplication_direct_73
-- reg_a = a3_X; reg_b = b3_X; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001110000000000100000100000011111001101100011",
--  (74) multiplication_direct_74
-- reg_a = a4_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000011111001010000011",
--  (75) multiplication_direct_75
-- reg_a = a2_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000011111010001000011",
--  (76) multiplication_direct_76
-- reg_a = a5_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000011111000110100011",
--  (77) multiplication_direct_77
-- reg_a = a1_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"001100100001110000000000100000000000011111010100100011",
--  (78) multiplication_direct_78
-- -- In case of size 7
-- reg_a = a6_X; reg_b = b0_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001110000000000100000000000111111000011000011",
--  (79) multiplication_direct_79
-- reg_a = a0_X; reg_b = b6_X; reg_acc = reg_o; o6_0 = reg_o; Enable sign b; operation : a*b + acc;
"000000100001110000010000100000000001011111011000000011",
--  (80) multiplication_direct_80
-- reg_a = a4_X; reg_b = b3_X; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001110000000000100000100000000011101110000011",
--  (81) multiplication_direct_81
-- reg_a = a3_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000011110001100011",
--  (82) multiplication_direct_82
-- reg_a = a5_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000011101010100011",
--  (83) multiplication_direct_83
-- reg_a = a2_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000011110101000011",
--  (84) multiplication_direct_84
-- reg_a = a6_X; reg_b = b1_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001110000000000100000000000100011100111000011",
--  (85) multiplication_direct_85
-- reg_a = a1_X; reg_b = b6_X; reg_acc = reg_o; o7_0 = reg_o; Enable sign b; operation : a*b + acc; Increment base address o;
"000000100001110010010000100000000001000011111000100011",
--  (86) multiplication_direct_86
-- reg_a = a4_X; reg_b = b4_X; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001110000000000100000100000000100010010000011",
--  (87) multiplication_direct_87
-- reg_a = a5_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001110100011",
--  (88) multiplication_direct_88
-- reg_a = a3_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010101100011",
--  (89) multiplication_direct_89
-- reg_a = a6_X; reg_b = b2_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001110000000000100000000000100100001011000011",
--  (90) multiplication_direct_90
-- reg_a = a2_X; reg_b = b6_X; reg_acc = reg_o; o8_0 = reg_o; Enable sign b; operation : a*b + acc;
"000000100001110000010000100000000001000100011001000011",
--  (91) multiplication_direct_91
-- reg_a = a5_X; reg_b = b4_X; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001110000000000100000100000001000110010100011",
--  (92) multiplication_direct_92
-- reg_a = a4_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000001000110110000011",
--  (93) multiplication_direct_93
-- reg_a = a6_X; reg_b = b3_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001110000000000100000000000101000101111000011",
--  (94) multiplication_direct_94
-- reg_a = a3_X; reg_b = b6_X; reg_acc = reg_o; o9_0 = reg_o; Enable sign b; operation : a*b + acc;
"000000100001110000010000100000000001001000111001100011",
--  (95) multiplication_direct_95
-- reg_a = a5_X; reg_b = b5_X; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001110000000000100000100000001101010110100011",
--  (96) multiplication_direct_96
-- reg_a = a6_X; reg_b = b4_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001110000000000100000000000101101010011000011",
--  (97) multiplication_direct_97
-- reg_a = a4_X; reg_b = b6_X; reg_acc = reg_o; o10_0 = reg_o; Enable sign b; operation : a*b + acc;
"000000100001110000010000100000000001001101011010000011",
--  (98) multiplication_direct_98
-- reg_a = a6_X; reg_b = b5_X; reg_acc = reg_o >> 256; Enable sign a; operation : a*b + acc;
"000000100001110000000000100000100000110001110111000011",
--  (99) multiplication_direct_99
-- reg_a = a5_X; reg_b = b6_X; reg_acc = reg_o; o11_0 = reg_o; Enable sign b; operation : a*b + acc;
"000000100001110000010000100000000001010001111010100011",
--  (100) multiplication_direct_100
-- reg_a = a6_X; reg_b = b6_X; reg_acc = reg_o >> 256; o12_X = reg_o; o13_X = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001110001110000100000100001110110011011000011",
--  (101) multiplication_direct_101
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (102) multiplication_direct_102
-- -- In case of size 8
-- reg_a = a6_X; reg_b = b0_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000011111000011000011",
--  (103) multiplication_direct_103
-- reg_a = a0_X; reg_b = b6_X; reg_acc = reg_o; o6_0 = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000011111011000000011",
--  (104) multiplication_direct_104
-- reg_a = a4_X; reg_b = b3_X; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001111000000000100000100000000011101110000011",
--  (105) multiplication_direct_105
-- reg_a = a3_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000011110001100011",
--  (106) multiplication_direct_106
-- reg_a = a5_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000011101010100011",
--  (107) multiplication_direct_107
-- reg_a = a2_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000011110101000011",
--  (108) multiplication_direct_108
-- reg_a = a6_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000011100111000011",
--  (109) multiplication_direct_109
-- reg_a = a1_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000011111000100011",
--  (110) multiplication_direct_110
-- reg_a = a7_X; reg_b = b0_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001111000000000100000000000100011100011100011",
--  (111) multiplication_direct_111
-- reg_a = a0_X; reg_b = b7_X; reg_acc = reg_o; o7_0 = reg_o; Enable sign b; operation : a*b + acc; Increment base address o;
"000000100001111010010000100000000001000011111100000011",
--  (112) multiplication_direct_112
-- reg_a = a4_X; reg_b = b4_X; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001111000000000100000100000000100010010000011",
--  (113) multiplication_direct_113
-- reg_a = a5_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001110100011",
--  (114) multiplication_direct_114
-- reg_a = a3_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010101100011",
--  (115) multiplication_direct_115
-- reg_a = a6_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001011000011",
--  (116) multiplication_direct_116
-- reg_a = a2_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011001000011",
--  (117) multiplication_direct_117
-- reg_a = a7_X; reg_b = b1_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001111000000000100000000000100100000111100011",
--  (118) multiplication_direct_118
-- reg_a = a1_X; reg_b = b7_X; reg_acc = reg_o; o8_0 = reg_o; Enable sign b; operation : a*b + acc;
"000000100001111000010000100000000001000100011100100011",
--  (119) multiplication_direct_119
-- reg_a = a5_X; reg_b = b4_X; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001111000000000100000100000001000110010100011",
--  (120) multiplication_direct_120
-- reg_a = a4_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000001000110110000011",
--  (121) multiplication_direct_121
-- reg_a = a6_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000001000101111000011",
--  (122) multiplication_direct_122
-- reg_a = a3_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000001000111001100011",
--  (123) multiplication_direct_123
-- reg_a = a7_X; reg_b = b2_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001111000000000100000000000101000101011100011",
--  (124) multiplication_direct_124
-- reg_a = a2_X; reg_b = b7_X; reg_acc = reg_o; o9_0 = reg_o; Enable sign b; operation : a*b + acc;
"000000100001111000010000100000000001001000111101000011",
--  (125) multiplication_direct_125
-- reg_a = a5_X; reg_b = b5_X; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001111000000000100000100000001101010110100011",
--  (126) multiplication_direct_126
-- reg_a = a6_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000001101010011000011",
--  (127) multiplication_direct_127
-- reg_a = a4_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000001101011010000011",
--  (128) multiplication_direct_128
-- reg_a = a7_X; reg_b = b3_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001111000000000100000000000101101001111100011",
--  (129) multiplication_direct_129
-- reg_a = a3_X; reg_b = b7_X; reg_acc = reg_o; o10_0 = reg_o; Enable sign b; operation : a*b + acc;
"000000100001111000010000100000000001001101011101100011",
--  (130) multiplication_direct_130
-- reg_a = a6_X; reg_b = b5_X; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001111000000000100000100000010001110111000011",
--  (131) multiplication_direct_131
-- reg_a = a5_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000010001111010100011",
--  (132) multiplication_direct_132
-- reg_a = a7_X; reg_b = b4_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001111000000000100000000000110001110011100011",
--  (133) multiplication_direct_133
-- reg_a = a4_X; reg_b = b7_X; reg_acc = reg_o; o11_0 = reg_o; Enable sign b; operation : a*b + acc;
"000000100001111000010000100000000001010001111110000011",
--  (134) multiplication_direct_134
-- reg_a = a6_X; reg_b = b6_X; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001111000000000100000100000010110011011000011",
--  (135) multiplication_direct_135
-- reg_a = a7_X; reg_b = b5_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001111000000000100000000000110110010111100011",
--  (136) multiplication_direct_136
-- reg_a = a5_X; reg_b = b7_X; reg_acc = reg_o; o12_0 = reg_o; Enable sign b; operation : a*b + acc;
"000000100001111000010000100000000001010110011110100011",
--  (137) multiplication_direct_137
-- reg_a = a7_X; reg_b = b6_X; reg_acc = reg_o >> 256; Enable sign a; operation : a*b + acc;
"000000100001111000000000100000100000111010111011100011",
--  (138) multiplication_direct_138
-- reg_a = a6_X; reg_b = b7_X; reg_acc = reg_o; o13_0 = reg_o; Enable sign b; operation : a*b + acc;
"000000100001111000010000100000000001011010111111000011",
--  (139) multiplication_direct_139
-- reg_a = a7_X; reg_b = b7_X; reg_acc = reg_o >> 256; o14_X = reg_o; o15_X = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001111001110000100000100001111111011111100011",
--  (140) multiplication_direct_140
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (141) square_direct_0
-- -- In case of size 1
-- reg_a = a0_X; reg_b = a0_X; reg_acc = 0; o0_X = reg_o; o1_X = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001000001110000100000010001100100000000000011",
--  (142) square_direct_1
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (143) square_direct_2
-- -- In case of sizes 2, 3, 4, 5, 6, 7, 8
-- reg_a = a0_X; reg_b = a0_X; reg_acc = 0; o0_X = reg_o; operation : a*b + acc;
"000010000001001000010000100000010000000100000000000011",
--  (144) square_direct_3
-- -- In case of size 2
-- reg_a = a1_X; reg_b = a0_X; reg_acc = reg_o >> 256; o1_X = reg_o; Enable sign a; operation : 2*a*b + acc;
"000000100001001000010100100000100000101000100000100011",
--  (145) square_direct_4
-- reg_a = a1_X; reg_b = a1_X; reg_acc = reg_o >> 256; o2_X = reg_o; o3_X = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001001001110000100000100001101101000100100011",
--  (146) square_direct_5
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (147) square_direct_6
-- -- Other cases
-- reg_a = a1_X; reg_b = a0_X; reg_acc = reg_o >> 256; o1_X = reg_o; operation : 2*a*b + acc;
"000000100001010000010100100000100000001000100000100011",
--  (148) square_direct_7
-- reg_a = a1_X; reg_b = a1_X; reg_acc = reg_o >> 256; operation : a*b + acc;
"000010100001010000000000100000100000001101000100100011",
--  (149) square_direct_8
-- -- In case of size 3
-- reg_a = a0_X; reg_b = a2_X; reg_acc = reg_o; o2_X = reg_o; Enable sign b; operation : 2*a*b + acc;
"000000100001010000010100100000000001001101001000000011",
--  (150) square_direct_9
-- reg_a = a2_X; reg_b = a1_X; reg_acc = reg_o >> 256; o3_X = reg_o; Enable sign a; operation : 2*a*b + acc;
"000000100001010000010100100000100000110001100101000011",
--  (151) square_direct_10
-- reg_a = a2_X; reg_b = a2_X; reg_acc = reg_o >> 256; o4_X = reg_o; o5_X = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001010001110000100000100001110110001001000011",
--  (152) square_direct_11
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (153) square_direct_12
-- -- Other cases
-- reg_a = a0_X; reg_b = a2_X; reg_acc = reg_o; o2_X = reg_o; operation : 2*a*b + acc;
"000000100001011000010100100000000000001101001000000011",
--  (154) square_direct_13
-- reg_a = a2_X; reg_b = a1_X; reg_acc = reg_o >> 256; operation : 2*a*b + acc;
"000011100001011000000100100000100000010001100101000011",
--  (155) square_direct_14
-- -- In case of size 4
-- reg_a = a3_X; reg_b = a0_X; reg_acc = reg_o; o3_X = reg_o; Enable sign a; operation : 2*a*b + acc;
"000000100001011000010100100000000000110001100001100011",
--  (156) square_direct_15
-- reg_a = a2_X; reg_b = a2_X; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001011000000000100000100000010110001001000011",
--  (157) square_direct_16
-- reg_a = a3_X; reg_b = a1_X; reg_acc = reg_o; o4_X = reg_o; Enable sign a; operation : 2*a*b + acc;
"000000100001011000010100100000000000110110000101100011",
--  (158) square_direct_17
-- reg_a = a3_X; reg_b = a2_X; reg_acc = reg_o >> 256; o5_X = reg_o; Enable sign a; operation : 2*a*b + acc;
"000000100001011000010100100000100000111010101001100011",
--  (159) square_direct_18
-- reg_a = a3_X; reg_b = a3_X; reg_acc = reg_o >> 256; o6_X = reg_o; o7_X = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001011001110000100000100001111111001101100011",
--  (160) square_direct_19
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (161) square_direct_20
-- -- Other cases
-- reg_a = a3_X; reg_b = a0_X; reg_acc = reg_o; o3_X = reg_o; operation : 2*a*b + acc;
"000000100001100000010100100000000000010001100001100011",
--  (162) square_direct_21
-- reg_a = a2_X; reg_b = a2_X; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001100000000000100000100000010110001001000011",
--  (163) square_direct_22
-- reg_a = a3_X; reg_b = a1_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000100100001100000000100100000000000010110000101100011",
--  (164) square_direct_23
-- -- In case of size 5
-- reg_a = a4_X; reg_b = a0_X; reg_acc = reg_o; o4_X = reg_o; Enable sign a; operation : 2*a*b + acc;
"000000100001100000010100100000000000110110000010000011",
--  (165) square_direct_24
-- reg_a = a3_X; reg_b = a2_X; reg_acc = reg_o >> 256; operation : 2*a*b + acc;
"000000100001100000000100100000100000011010101001100011",
--  (166) square_direct_25
-- reg_a = a4_X; reg_b = a1_X; reg_acc = reg_o; o5_X = reg_o; Enable sign a; operation : 2*a*b + acc;
"000000100001100000010100100000000000111010100110000011",
--  (167) square_direct_26
-- reg_a = a3_X; reg_b = a3_X; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001100000000000100000100000011111011011000011",
--  (168) square_direct_27
-- reg_a = a4_X; reg_b = a2_X; reg_acc = reg_o; o6_X = reg_o; Enable sign a; operation : 2*a*b + acc;
"000000100001100000010100100000000000111111001010000011",
--  (169) square_direct_28
-- reg_a = a4_X; reg_b = a3_X; reg_acc = reg_o >> 256; o7_X = reg_o; Enable sign a; operation : 2*a*b + acc; Increase base address o;
"000000100001100010010100100000100000100011101110000011",
--  (170) square_direct_29
-- reg_a = a4_X; reg_b = a4_X; reg_acc = reg_o >> 256; o8_X = reg_o; o9_X = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001100001110000100000100001100100010010000011",
--  (171) square_direct_30
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (172) square_direct_31
-- -- Other cases
-- reg_a = a4_X; reg_b = a0_X; reg_acc = reg_o; o4_X = reg_o; operation : 2*a*b + acc;
"000000100001101000010100100000000000010110000010000011",
--  (173) square_direct_32
-- reg_a = a3_X; reg_b = a2_X; reg_acc = reg_o >> 256; operation : 2*a*b + acc;
"000000100001101000000100100000100000010110001001100011",
--  (174) square_direct_33
-- reg_a = a4_X; reg_b = a1_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000110000001101000000100100000000000011010100110000011",
--  (175) square_direct_34
-- -- In case of size 6
-- reg_a = a5_X; reg_b = a0_X; reg_acc = reg_o; o5_X = reg_o; Enable sign a; operation : 2*a*b + acc;
"000000100001101000010100100000000000111010100010100011",
--  (176) square_direct_35
-- reg_a = a3_X; reg_b = a3_X; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001101000000000100000100000011111001101100011",
--  (177) square_direct_36
-- reg_a = a4_X; reg_b = a2_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001101000000100100000000000011111001010000011",
--  (178) square_direct_37
-- reg_a = a5_X; reg_b = a1_X; reg_acc = reg_o; o6_X = reg_o; Enable sign a; operation : 2*a*b + acc;
"000000100001101000010100100000000000111011000110100011",
--  (179) square_direct_38
-- reg_a = a4_X; reg_b = a3_X; reg_acc = reg_o >> 256; operation : 2*a*b + acc;
"000000100001101000000100100000100000000011101110000011",
--  (180) square_direct_39
-- reg_a = a5_X; reg_b = a2_X; reg_acc = reg_o; o7_X = reg_o; Enable sign a; operation : 2*a*b + acc; Increase base address o;
"000000100001101010010100100000000000100011101010100011",
--  (181) square_direct_40
-- reg_a = a4_X; reg_b = a4_X; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001101000000000100000100000000100010010000011",
--  (182) square_direct_41
-- reg_a = a5_X; reg_b = a3_X; reg_acc = reg_o; o8_X = reg_o; Enable sign a; operation : 2*a*b + acc;
"000000100001101000010100100000000000100100001110100011",
--  (183) square_direct_42
-- reg_a = a5_X; reg_b = a4_X; reg_acc = reg_o >> 256; o9_X = reg_o; Enable sign a; operation : 2*a*b + acc;
"000000100001101000010100100000100000101000110010100011",
--  (184) square_direct_43
-- reg_a = a5_X; reg_b = a5_X; reg_acc = reg_o >> 256; o10_X = reg_o; o11_X = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001101001110000100000100001101101010110100011",
--  (185) square_direct_44
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (186) square_direct_45
-- -- Other cases
-- reg_a = a5_X; reg_b = a0_X; reg_acc = reg_o; o5_X = reg_o; operation : 2*a*b + acc;
"000000100001110000010100100000000000011010100010100011",
--  (187) square_direct_46
-- reg_a = a3_X; reg_b = a3_X; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001110000000000100000100000011111001101100011",
--  (188) square_direct_47
-- reg_a = a4_X; reg_b = a2_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001110000000100100000000000011111001010000011",
--  (189) square_direct_48
-- reg_a = a5_X; reg_b = a1_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000111100001110000000100100000000000011111000110100011",
--  (190) square_direct_49
-- -- In case of size 7
-- reg_a = a6_X; reg_b = a0_X; reg_acc = reg_o; o6_X = reg_o; Enable sign a; operation : 2*a*b + acc;
"000000100001110000010100100000000000111111000011000011",
--  (191) square_direct_50
-- reg_a = a4_X; reg_b = a3_X; reg_acc = reg_o >> 256; operation : 2*a*b + acc;
"000000100001110000000100100000100000000011101110000011",
--  (192) square_direct_51
-- reg_a = a5_X; reg_b = a2_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001110000000100100000000000000011101010100011",
--  (193) square_direct_52
-- reg_a = a6_X; reg_b = a1_X; reg_acc = reg_o; o7_X = reg_o; Enable sign a; operation : 2*a*b + acc; Increase base address o;
"000000100001110010010100100000000000100011100111000011",
--  (194) square_direct_53
-- reg_a = a4_X; reg_b = a4_X; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001110000000000100000100000000100010010000011",
--  (195) square_direct_54
-- reg_a = a5_X; reg_b = a3_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001110000000100100000000000000100001110100011",
--  (196) square_direct_55
-- reg_a = a6_X; reg_b = a2_X; reg_acc = reg_o; o8_X = reg_o; Enable sign a; operation : 2*a*b + acc;
"000000100001110000010100100000000000100100001011000011",
--  (197) square_direct_56
-- reg_a = a5_X; reg_b = a4_X; reg_acc = reg_o >> 256; operation : 2*a*b + acc;
"000000100001110000000100100000100000001000110010100011",
--  (198) square_direct_57
-- reg_a = a6_X; reg_b = a3_X; reg_acc = reg_o; o9_X = reg_o; Enable sign a; operation : 2*a*b + acc;
"000000100001110000010100100000000000101000101111000011",
--  (199) square_direct_58
-- reg_a = a5_X; reg_b = a5_X; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001110000000000100000100000001101010110100011",
--  (200) square_direct_59
-- reg_a = a6_X; reg_b = a4_X; reg_acc = reg_o; o10_X = reg_o; Enable sign a; operation : 2*a*b + acc;
"000000100001110000010100100000000000101101010011000011",
--  (201) square_direct_60
-- reg_a = a6_X; reg_b = a5_X; reg_acc = reg_o >> 256; o11_X = reg_o; Enable sign a; operation : 2*a*b + acc;
"000000100001110000010100100000100000110001110111000011",
--  (202) square_direct_61
-- reg_a = a6_X; reg_b = a6_X; reg_acc = reg_o >> 256; o12_X = reg_o; o13_X = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001110001110000100000100001110110011011000011",
--  (203) square_direct_62
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (204) square_direct_63
-- -- In case of size 8
-- reg_a = a6_X; reg_b = a0_X; reg_acc = reg_o; o6_X = reg_o; operation : 2*a*b + acc;
"000000100001111000010100100000000000011111000011000011",
--  (205) square_direct_64
-- reg_a = a4_X; reg_b = a3_X; reg_acc = reg_o >> 256; operation : 2*a*b + acc;
"000000100001111000000100100000100000000011101110000011",
--  (206) square_direct_65
-- reg_a = a5_X; reg_b = a2_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001111000000100100000000000000011101010100011",
--  (207) square_direct_66
-- reg_a = a6_X; reg_b = a1_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001111000000100100000000000000011100111000011",
--  (208) square_direct_67
-- reg_a = a7_X; reg_b = a0_X; reg_acc = reg_o; o7_X = reg_o; Enable sign a; operation : 2*a*b + acc; Increase base address o;
"000000100001111010010100100000000000100011100011100011",
--  (209) square_direct_68
-- reg_a = a4_X; reg_b = a4_X; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001111000000000100000100000000100010010000011",
--  (210) square_direct_69
-- reg_a = a5_X; reg_b = a3_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001111000000100100000000000000100001110100011",
--  (211) square_direct_70
-- reg_a = a6_X; reg_b = a2_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001111000000100100000000000000100001011000011",
--  (212) square_direct_71
-- reg_a = a7_X; reg_b = a1_X; reg_acc = reg_o; o8_X = reg_o; Enable sign a; operation : 2*a*b + acc;
"000000100001111000010100100000000000100100000111100011",
--  (213) square_direct_72
-- reg_a = a5_X; reg_b = a4_X; reg_acc = reg_o >> 256; operation : 2*a*b + acc;
"000000100001111000000100100000100000001000110010100011",
--  (214) square_direct_73
-- reg_a = a6_X; reg_b = a3_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001111000000100100000000000001000101111000011",
--  (215) square_direct_74
-- reg_a = a7_X; reg_b = a2_X; reg_acc = reg_o; o9_X = reg_o; Enable sign a; operation : 2*a*b + acc;
"000000100001111000010100100000000000101000101011100011",
--  (216) square_direct_75
-- reg_a = a5_X; reg_b = a5_X; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001111000000000100000100000001101010110100011",
--  (217) square_direct_76
-- reg_a = a6_X; reg_b = a4_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001111000000100100000000000001101010011000011",
--  (218) square_direct_77
-- reg_a = a7_X; reg_b = a3_X; reg_acc = reg_o; o10_X = reg_o; Enable sign a; operation : 2*a*b + acc;
"000000100001111000010100100000000000101101001111100011",
--  (219) square_direct_78
-- reg_a = a6_X; reg_b = a5_X; reg_acc = reg_o >> 256; operation : 2*a*b + acc;
"000000100001111000000100100000100000010001110111000011",
--  (220) square_direct_79
-- reg_a = a7_X; reg_b = a4_X; reg_acc = reg_o; o11_X = reg_o; Enable sign a; operation : 2*a*b + acc;
"000000100001111000010100100000000000110001110011100011",
--  (221) square_direct_80
-- reg_a = a6_X; reg_b = a6_X; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001111000000000100000100000010110011011000011",
--  (222) square_direct_81
-- reg_a = a7_X; reg_b = a5_X; reg_acc = reg_o; o12_X = reg_o; Enable sign a; operation : 2*a*b + acc;
"000000100001111000010100100000000000110110010111100011",
--  (223) square_direct_82
-- reg_a = a7_X; reg_b = a6_X; reg_acc = reg_o >> 256; o13_X = reg_o; Enable sign a; operation : 2*a*b + acc;
"000000100001111000010100100000100000111010111011100011",
--  (224) square_direct_83
-- reg_a = a7_X; reg_b = a7_X; reg_acc = reg_o >> 256; o14_X = reg_o; o15_X = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001111001110000100000100001111111011111100011",
--  (225) square_direct_84
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (226) multiplication_with_reduction_0
-- -- In case of size 1
-- reg_a = a0_X; reg_b = b0_X; reg_acc = 0; Enable sign a,b; operation : a*b + acc;
"000000100001000000000000100000010001100100000000000011",
--  (227) multiplication_with_reduction_1
-- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o0_X = reg_y; operation : keep accumulator;
"000000100001000000011000110000000100000100000000011011",
--  (228) multiplication_with_reduction_2
-- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
"000000100001000000000000100000000010000100000000010011",
--  (229) multiplication_with_reduction_3
-- reg_a = 0; reg_b = 0; reg_acc = reg_o >> 256; o0_X = reg_o; operation : a*b + acc;
"000000100001000000010000100000101110000100000000000011",
--  (230) multiplication_with_reduction_4
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (231) multiplication_with_reduction_5
-- -- In case of sizes 2, 3, 4, 5, 6, 7, 8
-- reg_a = a0_X; reg_b = b0_X; reg_acc = 0; operation : a*b + acc;
"000000100001001000000000100000010000000100000000000011",
--  (232) multiplication_with_reduction_6
-- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o0_X = reg_y; operation : keep accumulator;
"000000100001001000011000110000000100000100000000011011",
--  (233) multiplication_with_reduction_7
-- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
"000000100001001000000000100000000010000100000000010011",
--  (234) multiplication_with_reduction_8
--reg_a = o0_X; reg_b = prime1; reg_acc = reg_o >> 256; operation : a*b + acc;
"000100000001001000000000100000100000000100000100010111",
--  (235) multiplication_with_reduction_9
-- -- In case of size 2
-- reg_a = a0_X; reg_b = b1_X; reg_acc = reg_o; Enable sign b; operation : a*b + acc;
"000000100001001000000000100000000001000100000100000011",
--  (236) multiplication_with_reduction_10
-- reg_a = a1_X; reg_b = b0_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001001000000000100000000000100100000000100011",
--  (237) multiplication_with_reduction_11
-- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o1_X = reg_y; operation : keep accumulator;
"000000100001001000011000110000000100001000100000011011",
--  (238) multiplication_with_reduction_12
-- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
"000000100001001000000000100000000010000100000000010011",
--  (239) multiplication_with_reduction_13
-- reg_a = a1_X; reg_b = b1_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001001000000000100000100001100100000100100011",
--  (240) multiplication_with_reduction_14
-- reg_a = o1_X; reg_b = prime1; reg_acc = reg_o; o0_X = reg_o; o1_X = reg_o >> 256; operation : a*b + acc;
"000000100001001001110000100000000000000100000100110111",
--  (241) multiplication_with_reduction_15
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (242) multiplication_with_reduction_16
-- -- Other cases
-- reg_a = a0_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001010000000000100000000000000100000100000011",
--  (243) multiplication_with_reduction_17
-- reg_a = a1_X; reg_b = b0_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001010000000000100000000000000100000000100011",
--  (244) multiplication_with_reduction_18
-- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o1_X = reg_y; operation : keep accumulator;
"000000100001010000011000110000000100001000100000011011",
--  (245) multiplication_with_reduction_19
-- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
"000000100001010000000000100000000010000100000000010011",
--  (246) multiplication_with_reduction_20
-- reg_a = o0_X; reg_b = prime2; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001010000000000100000100000000100001000010111",
--  (247) multiplication_with_reduction_21
-- reg_a = a1_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001010000000000100000000000000100000100100011",
--  (248) multiplication_with_reduction_22
-- reg_a = o1_X; reg_b = prime1; reg_acc = reg_o; operation : a*b + acc;
"000110000001010000000000100000000000000100000100110111",
--  (249) multiplication_with_reduction_23
-- -- In case of size 3
-- reg_a = a0_X; reg_b = b2_X; reg_acc = reg_o; Enable sign b; operation : a*b + acc;
"000000100001010000000000100000000001000100001000000011",
--  (250) multiplication_with_reduction_24
-- reg_a = a2_X; reg_b = b0_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001010000000000100000000000100100000001000011",
--  (251) multiplication_with_reduction_25
-- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o2_X = reg_y; operation : keep accumulator;
"000000100001010000011000110000000100001101000000011011",
--  (252) multiplication_with_reduction_26
-- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
"000000100001010000000000100000000010000100000000010011",
--  (253) multiplication_with_reduction_27
-- reg_a = a1_X; reg_b = b2_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001010000000000100000100001000100001000100011",
--  (254) multiplication_with_reduction_28
-- reg_a = o1_X; reg_b = prime2; reg_acc = reg_o; operation : a*b + acc;
"000000100001010000000000100000000000000100001000110111",
--  (255) multiplication_with_reduction_29
-- reg_a = a2_X; reg_b = b1_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001010000000000100000000000100100000101000011",
--  (256) multiplication_with_reduction_30
-- reg_a = o2_X; reg_b = prime1; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
"000000100001010000010000100000000000000100000101010111",
--  (257) multiplication_with_reduction_31
-- reg_a = a2_X; reg_b = b2_X; reg_acc = reg_o >> 256; Enable sign a, b; operation : a*b + acc;
"000000100001010000000000100000100001100100001001000011",
--  (258) multiplication_with_reduction_32
-- reg_a = o2_X; reg_b = prime2; reg_acc = reg_o; o1_X = reg_o; o2_X = reg_o >> 256; operation : a*b + acc;
"000000100001010001110000100000000000001000101001010111",
--  (259) multiplication_with_reduction_33
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (260) multiplication_with_reduction_34
-- -- Other cases
-- reg_a = a0_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001011000000000100000000000000100001000000011",
--  (261) multiplication_with_reduction_35
-- reg_a = a2_X; reg_b = b0_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001011000000000100000000000000100000001000011",
--  (262) multiplication_with_reduction_36
-- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o2_X = reg_y; operation : keep accumulator;
"000000100001011000011000110000000100001101000000011011",
--  (263) multiplication_with_reduction_37
-- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
"000000100001011000000000100000000010000100000000010011",
--  (264) multiplication_with_reduction_38
-- reg_a = o0_X; reg_b = prime3; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001011000000000100000100000000100001100010111",
--  (265) multiplication_with_reduction_39
-- reg_a = a1_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001011000000000100000000000000100001000100011",
--  (266) multiplication_with_reduction_40
-- reg_a = o1_X; reg_b = prime2; reg_acc = reg_o; operation : a*b + acc;
"000000100001011000000000100000000000000100001000110111",
--  (267) multiplication_with_reduction_41
-- reg_a = a2_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001011000000000100000000000000100000101000011",
--  (268) multiplication_with_reduction_42
-- reg_a = o2_X; reg_b = prime1; reg_acc = reg_o; operation : a*b + acc;
"001001000001011000000000100000000000000100000101010111",
--  (269) multiplication_with_reduction_43
-- -- In case of size 4
-- reg_a = a0_X; reg_b = b3_X; reg_acc = reg_o; Enable sign b; operation : a*b + acc;
"000000100001011000000000100000000001000100001100000011",
--  (270) multiplication_with_reduction_44
-- reg_a = a3_X; reg_b = b0_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001011000000000100000000000100100000001100011",
--  (271) multiplication_with_reduction_45
-- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o3_X = reg_y; operation : keep accumulator;
"000000100001011000011000110000000100000001100000011011",
--  (272) multiplication_with_reduction_46
-- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
"000000100001011000000000100000000010000100000000010011",
--  (273) multiplication_with_reduction_47
-- reg_a = a1_X; reg_b = b3_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001011000000000100000100001000100001100100011",
--  (274) multiplication_with_reduction_48
-- reg_a = o1_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
"000000100001011000000000100000000000000100001100110111",
--  (275) multiplication_with_reduction_49
-- reg_a = a2_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001011000000000100000000000000100001001000011",
--  (276) multiplication_with_reduction_50
-- reg_a = o2_X; reg_b = prime2; reg_acc = reg_o; operation : a*b + acc;
"000000100001011000000000100000000000000100001001010111",
--  (277) multiplication_with_reduction_51
-- reg_a = a3_X; reg_b = b1_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001011000000000100000000000100100000101100011",
--  (278) multiplication_with_reduction_52
-- reg_a = o3_X; reg_b = prime1; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
"000000100001011000010000100000000000000100000101110111",
--  (279) multiplication_with_reduction_53
-- reg_a = a2_X; reg_b = b3_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001011000000000100000100001000100001101000011",
--  (280) multiplication_with_reduction_54
-- reg_a = o2_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
"000000100001011000000000100000000000000100001101010111",
--  (281) multiplication_with_reduction_55
-- reg_a = a3_X; reg_b = b2_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001011000000000100000000000100100001001100011",
--  (282) multiplication_with_reduction_56
-- reg_a = o3_X; reg_b = prime2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
"000000100001011000010000100000000000001000101001110111",
--  (283) multiplication_with_reduction_57
-- reg_a = a3_X; reg_b = b3_X; reg_acc = reg_o >> 256; Enable sign a, b; operation : a*b + acc;
"000000100001011000000000100000100001100100001101100011",
--  (284) multiplication_with_reduction_58
-- reg_a = o3_X; reg_b = prime3; reg_acc = reg_o; o2_X = reg_o; o3_0 = reg_o >> 256; operation : a*b + acc;
"000000100001011001110000100000000000001101001101110111",
--  (285) multiplication_with_reduction_59
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (286) multiplication_with_reduction_60
-- -- Other cases
-- reg_a = a0_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001100000011",
--  (287) multiplication_with_reduction_61
-- reg_a = a3_X; reg_b = b0_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100000001100011",
--  (288) multiplication_with_reduction_62
-- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o3_X = reg_y; operation : keep accumulator;
"000000100001100000011000110000000100010001100000011011",
--  (289) multiplication_with_reduction_63
-- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000010000100000000010011",
--  (290) multiplication_with_reduction_64
-- reg_a = o0_X; reg_b = prime4; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001100000000000100000100000000100010000010111",
--  (291) multiplication_with_reduction_65
-- reg_a = a1_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001100100011",
--  (292) multiplication_with_reduction_66
-- reg_a = o1_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001100110111",
--  (293) multiplication_with_reduction_67
-- reg_a = a2_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001001000011",
--  (294) multiplication_with_reduction_68
-- reg_a = o2_X; reg_b = prime2; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001001010111",
--  (295) multiplication_with_reduction_69
-- reg_a = a3_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100000101100011",
--  (296) multiplication_with_reduction_70
-- reg_a = o3_X; reg_b = prime1; reg_acc = reg_o; operation : a*b + acc;
"001101000001100000000000100000000000000100000101110111",
--  (297) multiplication_with_reduction_71
-- -- In case of size 5
-- reg_a = a0_X; reg_b = b4_X; reg_acc = reg_o; Enable sign b; operation : a*b + acc;
"000000100001100000000000100000000001000100010000000011",
--  (298) multiplication_with_reduction_72
-- reg_a = a4_X; reg_b = b0_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001100000000000100000000000100100000010000011",
--  (299) multiplication_with_reduction_73
-- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o4_X = reg_y; operation : keep accumulator;
"000000100001100000011000110000000100010110000000011011",
--  (300) multiplication_with_reduction_74
-- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000010000100000000010011",
--  (301) multiplication_with_reduction_75
-- reg_a = a1_X; reg_b = b4_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001100000000000100000100001000100010000100011",
--  (302) multiplication_with_reduction_76
-- reg_a = o1_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100010000110111",
--  (303) multiplication_with_reduction_77
-- reg_a = a2_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001101000011",
--  (304) multiplication_with_reduction_78
-- reg_a = o2_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001101010111",
--  (305) multiplication_with_reduction_79
-- reg_a = a3_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001001100011",
--  (306) multiplication_with_reduction_80
-- reg_a = o3_X; reg_b = prime2; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001001110111",
--  (307) multiplication_with_reduction_81
-- reg_a = a4_X; reg_b = b1_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001100000000000100000000000100100000110000011",
--  (308) multiplication_with_reduction_82
-- reg_a = o4_X; reg_b = prime1; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
"000000100001100000010000100000000000000100000110010111",
--  (309) multiplication_with_reduction_83
-- reg_a = a2_X; reg_b = b4_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001100000000000100000100001000100010001000011",
--  (310) multiplication_with_reduction_84
-- reg_a = o2_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100010001010111",
--  (311) multiplication_with_reduction_85
-- reg_a = a3_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001101100011",
--  (312) multiplication_with_reduction_86
-- reg_a = o3_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001101110111",
--  (313) multiplication_with_reduction_87
-- reg_a = a4_X; reg_b = b2_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001100000000000100000000000100100001010000011",
--  (314) multiplication_with_reduction_88
-- reg_a = o4_X; reg_b = prime2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
"000000100001100000010000100000000000001000101010010111",
--  (315) multiplication_with_reduction_89
-- reg_a = a3_X; reg_b = b4_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001100000000000100000100001000100010001100011",
--  (316) multiplication_with_reduction_90
-- reg_a = o3_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100010001110111",
--  (317) multiplication_with_reduction_91
-- reg_a = a4_X; reg_b = b3_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001100000000000100000000000100100001110000011",
--  (318) multiplication_with_reduction_92
-- reg_a = o4_X; reg_b = prime3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
"000000100001100000010000100000000000001101001110010111",
--  (319) multiplication_with_reduction_93
-- reg_a = a4_X; reg_b = b4_X; reg_acc = reg_o >> 256; Enable sign a, b; operation : a*b + acc;
"000000100001100000000000100000100001100100010010000011",
--  (320) multiplication_with_reduction_94
-- reg_a = o4_X; reg_b = prime4; reg_acc = reg_o; o3_X = reg_o; o4_0 = reg_o >> 256; operation : a*b + acc;
"000000100001100001110000100000000000010001110010010111",
--  (321) multiplication_with_reduction_95
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (322) multiplication_with_reduction_96
-- -- Other cases
-- reg_a = a0_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010000000011",
--  (323) multiplication_with_reduction_97
-- reg_a = a4_X; reg_b = b0_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100000010000011",
--  (324) multiplication_with_reduction_98
-- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o4_X = reg_y; operation : keep accumulator;
"000000100001101000011000110000000100010110000000011011",
--  (325) multiplication_with_reduction_99
-- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000010000100000000010011",
--  (326) multiplication_with_reduction_100
-- reg_a = o0_X; reg_b = prime5; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001101000000000100000100000000100010100010111",
--  (327) multiplication_with_reduction_101
-- reg_a = a1_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010000100011",
--  (328) multiplication_with_reduction_102
-- reg_a = o1_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010000110111",
--  (329) multiplication_with_reduction_103
-- reg_a = a2_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001101000011",
--  (330) multiplication_with_reduction_104
-- reg_a = o2_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001101010111",
--  (331) multiplication_with_reduction_105
-- reg_a = a3_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001001100011",
--  (332) multiplication_with_reduction_106
-- reg_a = o3_X; reg_b = prime2; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001001110111",
--  (333) multiplication_with_reduction_107
-- reg_a = a4_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100000110000011",
--  (334) multiplication_with_reduction_108
-- reg_a = o4_X; reg_b = prime1; reg_acc = reg_o; operation : a*b + acc;
"010010000001101000000000100000000000000100000110010111",
--  (335) multiplication_with_reduction_109
-- -- In case of size 6
-- reg_a = a0_X; reg_b = b5_X; reg_acc = reg_o; Enable sign b; operation : a*b + acc;
"000000100001101000000000100000000001000100010100000011",
--  (336) multiplication_with_reduction_110
-- reg_a = a5_X; reg_b = b0_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001101000000000100000000000100100000010100011",
--  (337) multiplication_with_reduction_111
-- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o5_X = reg_y; operation : keep accumulator;
"000000100001101000011000110000000100011010100000011011",
--  (338) multiplication_with_reduction_112
-- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000010000100000000010011",
--  (339) multiplication_with_reduction_113
-- reg_a = a1_X; reg_b = b5_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001101000000000100000100001000100010100100011",
--  (340) multiplication_with_reduction_114
-- reg_a = o1_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010100110111",
--  (341) multiplication_with_reduction_115
-- reg_a = a2_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010001000011",
--  (342) multiplication_with_reduction_116
-- reg_a = o2_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010001010111",
--  (343) multiplication_with_reduction_117
-- reg_a = a3_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001101100011",
--  (344) multiplication_with_reduction_118
-- reg_a = o3_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001101110111",
--  (345) multiplication_with_reduction_119
-- reg_a = a4_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001010000011",
--  (346) multiplication_with_reduction_120
-- reg_a = o4_X; reg_b = prime2; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001010010111",
--  (347) multiplication_with_reduction_121
-- reg_a = a5_X; reg_b = b1_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001101000000000100000000000100100000110100011",
--  (348) multiplication_with_reduction_122
-- reg_a = o5_X; reg_b = prime1; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
"000000100001101000010000100000000000000100000110110111",
--  (349) multiplication_with_reduction_123
-- reg_a = a2_X; reg_b = b5_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001101000000000100000100001000100010101000011",
--  (350) multiplication_with_reduction_124
-- reg_a = o2_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010101010111",
--  (351) multiplication_with_reduction_125
-- reg_a = a3_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010001100011",
--  (352) multiplication_with_reduction_126
-- reg_a = o3_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010001110111",
--  (353) multiplication_with_reduction_127
-- reg_a = a4_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001110000011",
--  (354) multiplication_with_reduction_128
-- reg_a = o4_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001110010111",
--  (355) multiplication_with_reduction_129
-- reg_a = a5_X; reg_b = b2_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001101000000000100000000000100100001010100011",
--  (356) multiplication_with_reduction_130
-- reg_a = o5_X; reg_b = prime2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
"000000100001101000010000100000000000001000101010110111",
--  (357) multiplication_with_reduction_131
-- reg_a = a3_X; reg_b = b5_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001101000000000100000100001000100010101100011",
--  (358) multiplication_with_reduction_132
-- reg_a = o3_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010101110111",
--  (359) multiplication_with_reduction_133
-- reg_a = a4_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010010000011",
--  (360) multiplication_with_reduction_134
-- reg_a = o4_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010010010111",
--  (361) multiplication_with_reduction_135
-- reg_a = a5_X; reg_b = b3_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001101000000000100000000000100100001110100011",
--  (362) multiplication_with_reduction_136
-- reg_a = o5_X; reg_b = prime3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
"000000100001101000010000100000000000001101001110110111",
--  (363) multiplication_with_reduction_137
-- reg_a = a4_X; reg_b = b5_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001101000000000100000100001000100010110000011",
--  (364) multiplication_with_reduction_138
-- reg_a = o4_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010110010111",
--  (365) multiplication_with_reduction_139
-- reg_a = a5_X; reg_b = b4_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001101000000000100000000000100100010010100011",
--  (366) multiplication_with_reduction_140
-- reg_a = o5_X; reg_b = prime4; reg_acc = reg_o; o3_X = reg_o; operation : a*b + acc;
"000000100001101000010000100000000000010001110010110111",
--  (367) multiplication_with_reduction_141
-- reg_a = a5_X; reg_b = b5_X; reg_acc = reg_o >> 256; Enable sign a, b; operation : a*b + acc;
"000000100001101000000000100000100001100100010110100011",
--  (368) multiplication_with_reduction_142
-- reg_a = o5_X; reg_b = prime5; reg_acc = reg_o; o4_X = reg_o; o5_0 = reg_o >> 256; operation : a*b + acc;
"000000100001101001110000100000000000010110010110110111",
--  (369) multiplication_with_reduction_143
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (370) multiplication_with_reduction_144
-- -- Other cases
-- reg_a = a0_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010100000011",
--  (371) multiplication_with_reduction_145
-- reg_a = a5_X; reg_b = b0_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100000010100011",
--  (372) multiplication_with_reduction_146
-- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o5_X = reg_y; operation : keep accumulator;
"000000100001110000011000110000000100011010100000011011",
--  (373) multiplication_with_reduction_147
-- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000010000100000000010011",
--  (374) multiplication_with_reduction_148
-- reg_a = o0_X; reg_b = prime6; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001110000000000100000100000000100011000010111",
--  (375) multiplication_with_reduction_149
-- reg_a = a1_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010100100011",
--  (376) multiplication_with_reduction_150
-- reg_a = o1_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010100110111",
--  (377) multiplication_with_reduction_151
-- reg_a = a2_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010001000011",
--  (378) multiplication_with_reduction_152
-- reg_a = o2_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010001010111",
--  (379) multiplication_with_reduction_153
-- reg_a = a3_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001101100011",
--  (380) multiplication_with_reduction_154
-- reg_a = o3_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001101110111",
--  (381) multiplication_with_reduction_155
-- reg_a = a4_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001010000011",
--  (382) multiplication_with_reduction_156
-- reg_a = o4_X; reg_b = prime2; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001010010111",
--  (383) multiplication_with_reduction_157
-- reg_a = a5_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100000110100011",
--  (384) multiplication_with_reduction_158
-- reg_a = o5_X; reg_b = prime1; reg_acc = reg_o; operation : a*b + acc;
"011000000001110000000000100000000000000100000110110111",
--  (385) multiplication_with_reduction_159
-- -- In case of size 7
-- reg_a = a0_X; reg_b = b6_X; reg_acc = reg_o; Enable sign b; operation : a*b + acc;
"000000100001110000000000100000000001000100011000000011",
--  (386) multiplication_with_reduction_160
-- reg_a = a6_X; reg_b = b0_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001110000000000100000000000100100000011000011",
--  (387) multiplication_with_reduction_161
-- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o6_X = reg_y; operation : keep accumulator;
"000000100001110000011000110000000100011111000000011011",
--  (388) multiplication_with_reduction_162
-- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000010000100000000010011",
--  (389) multiplication_with_reduction_163
-- reg_a = a1_X; reg_b = b6_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001110000000000100000100001000100011000100011",
--  (390) multiplication_with_reduction_164
-- reg_a = o1_X; reg_b = prime6; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100011000110111",
--  (391) multiplication_with_reduction_165
-- reg_a = a2_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010101000011",
--  (392) multiplication_with_reduction_166
-- reg_a = o2_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010101010111",
--  (393) multiplication_with_reduction_167
-- reg_a = a3_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010001100011",
--  (394) multiplication_with_reduction_168
-- reg_a = o3_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010001110111",
--  (395) multiplication_with_reduction_169
-- reg_a = a4_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001110000011",
--  (396) multiplication_with_reduction_170
-- reg_a = o4_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001110010111",
--  (397) multiplication_with_reduction_171
-- reg_a = a5_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001010100011",
--  (398) multiplication_with_reduction_172
-- reg_a = o5_X; reg_b = prime2; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001010110111",
--  (399) multiplication_with_reduction_173
-- reg_a = a6_X; reg_b = b1_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001110000000000100000000000100100000111000011",
--  (400) multiplication_with_reduction_174
-- reg_a = o6_X; reg_b = prime1; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
"000000100001110000010000100000000000000100000111010111",
--  (401) multiplication_with_reduction_175
-- reg_a = a2_X; reg_b = b6_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001110000000000100000100001000100011001000011",
--  (402) multiplication_with_reduction_176
-- reg_a = o2_X; reg_b = prime6; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100011001010111",
--  (403) multiplication_with_reduction_177
-- reg_a = a3_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010101100011",
--  (404) multiplication_with_reduction_178
-- reg_a = o3_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010101110111",
--  (405) multiplication_with_reduction_179
-- reg_a = a4_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010010000011",
--  (406) multiplication_with_reduction_180
-- reg_a = o4_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010010010111",
--  (407) multiplication_with_reduction_181
-- reg_a = a5_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001110100011",
--  (408) multiplication_with_reduction_182
-- reg_a = o5_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001110110111",
--  (409) multiplication_with_reduction_183
-- reg_a = a6_X; reg_b = b2_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001110000000000100000000000100100001011000011",
--  (410) multiplication_with_reduction_184
-- reg_a = o6_X; reg_b = prime2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
"000000100001110000010000100000000000001000101011010111",
--  (411) multiplication_with_reduction_185
-- reg_a = a3_X; reg_b = b6_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001110000000000100000100001000100011001100011",
--  (412) multiplication_with_reduction_186
-- reg_a = o3_X; reg_b = prime6; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100011001110111",
--  (413) multiplication_with_reduction_187
-- reg_a = a4_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010110000011",
--  (414) multiplication_with_reduction_188
-- reg_a = o4_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010110010111",
--  (415) multiplication_with_reduction_189
-- reg_a = a5_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010010100011",
--  (416) multiplication_with_reduction_190
-- reg_a = o5_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010010110111",
--  (417) multiplication_with_reduction_191
-- reg_a = a6_X; reg_b = b3_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001110000000000100000000000100100001111000011",
--  (418) multiplication_with_reduction_192
-- reg_a = o6_X; reg_b = prime3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
"000000100001110000010000100000000000001101001111010111",
--  (419) multiplication_with_reduction_193
-- reg_a = a4_X; reg_b = b6_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001110000000000100000100001000100011010000011",
--  (420) multiplication_with_reduction_194
-- reg_a = o4_X; reg_b = prime6; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100011010010111",
--  (421) multiplication_with_reduction_195
-- reg_a = a5_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010110100011",
--  (422) multiplication_with_reduction_196
-- reg_a = o5_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010110110111",
--  (423) multiplication_with_reduction_197
-- reg_a = a6_X; reg_b = b4_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001110000000000100000000000100100010011000011",
--  (424) multiplication_with_reduction_198
-- reg_a = o6_X; reg_b = prime4; reg_acc = reg_o; o3_X = reg_o; operation : a*b + acc;
"000000100001110000010000100000000000010001110011010111",
--  (425) multiplication_with_reduction_199
-- reg_a = a5_X; reg_b = b6_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001110000000000100000100001000100011010100011",
--  (426) multiplication_with_reduction_200
-- reg_a = o5_X; reg_b = prime6; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100011010110111",
--  (427) multiplication_with_reduction_201
-- reg_a = a6_X; reg_b = b5_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001110000000000100000000000100100010111000011",
--  (428) multiplication_with_reduction_202
-- reg_a = o6_X; reg_b = prime5; reg_acc = reg_o; o4_X = reg_o; operation : a*b + acc;
"000000100001110000010000100000000000010110010111010111",
--  (429) multiplication_with_reduction_203
-- reg_a = a6_X; reg_b = b6_X; reg_acc = reg_o >> 256; Enable sign a, b; operation : a*b + acc;
"000000100001110000000000100000100001100100011011000011",
--  (430) multiplication_with_reduction_204
-- reg_a = o6_X; reg_b = prime6; reg_acc = reg_o; o5_X = reg_o; o6_0 = reg_o >> 256; operation : a*b + acc;
"000000100001110001110000100000000000011010111011010111",
--  (431) multiplication_with_reduction_205
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (432) multiplication_with_reduction_206
-- -- In case of size 8
-- reg_a = a0_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011000000011",
--  (433) multiplication_with_reduction_207
-- reg_a = a6_X; reg_b = b0_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100000011000011",
--  (434) multiplication_with_reduction_208
-- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o6_X = reg_y; operation : keep accumulator;
"000000100001111000011000110000000100011111000000011011",
--  (435) multiplication_with_reduction_209
-- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000010000100000000010011",
--  (436) multiplication_with_reduction_210
-- reg_a = o0_X; reg_b = prime7; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001111000000000100000100000000100011100010111",
--  (437) multiplication_with_reduction_211
-- reg_a = a1_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011000100011",
--  (438) multiplication_with_reduction_212
-- reg_a = o1_X; reg_b = prime6; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011000110111",
--  (439) multiplication_with_reduction_213
-- reg_a = a2_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010101000011",
--  (440) multiplication_with_reduction_214
-- reg_a = o2_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010101010111",
--  (441) multiplication_with_reduction_215
-- reg_a = a3_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010001100011",
--  (442) multiplication_with_reduction_216
-- reg_a = o3_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010001110111",
--  (443) multiplication_with_reduction_217
-- reg_a = a4_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001110000011",
--  (444) multiplication_with_reduction_218
-- reg_a = o4_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001110010111",
--  (445) multiplication_with_reduction_219
-- reg_a = a5_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001010100011",
--  (446) multiplication_with_reduction_220
-- reg_a = o5_X; reg_b = prime2; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001010110111",
--  (447) multiplication_with_reduction_221
-- reg_a = a6_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100000111000011",
--  (448) multiplication_with_reduction_222
-- reg_a = o6_X; reg_b = prime1; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100000111010111",
--  (449) multiplication_with_reduction_223
-- reg_a = a0_X; reg_b = b7_X; reg_acc = reg_o; Enable sign b; operation : a*b + acc;
"000000100001111000000000100000000001000100011100000011",
--  (450) multiplication_with_reduction_224
-- reg_a = a7_X; reg_b = b0_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001111000000000100000000000100100000011100011",
--  (451) multiplication_with_reduction_225
-- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o7_X = reg_y; operation : keep accumulator;
"000000100001111000011000110000000100011111100000011011",
--  (452) multiplication_with_reduction_226
-- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000010000100000000010011",
--  (453) multiplication_with_reduction_227
-- reg_a = a1_X; reg_b = b7_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001111000000000100000100001000100011100100011",
--  (454) multiplication_with_reduction_228
-- reg_a = o1_X; reg_b = prime7; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011100110111",
--  (455) multiplication_with_reduction_229
-- reg_a = a2_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011001000011",
--  (456) multiplication_with_reduction_230
-- reg_a = o2_X; reg_b = prime6; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011001010111",
--  (457) multiplication_with_reduction_231
-- reg_a = a3_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010101100011",
--  (458) multiplication_with_reduction_232
-- reg_a = o3_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010101110111",
--  (459) multiplication_with_reduction_233
-- reg_a = a4_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010010000011",
--  (460) multiplication_with_reduction_234
-- reg_a = o4_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010010010111",
--  (461) multiplication_with_reduction_235
-- reg_a = a5_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001110100011",
--  (462) multiplication_with_reduction_236
-- reg_a = o5_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001110110111",
--  (463) multiplication_with_reduction_237
-- reg_a = a6_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001011000011",
--  (464) multiplication_with_reduction_238
-- reg_a = o6_X; reg_b = prime2; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001011010111",
--  (465) multiplication_with_reduction_239
-- reg_a = a7_X; reg_b = b1_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001111000000000100000000000100100000111100011",
--  (466) multiplication_with_reduction_240
-- reg_a = o7_X; reg_b = prime1; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000000100000111110111",
--  (467) multiplication_with_reduction_241
-- reg_a = a2_X; reg_b = b7_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001111000000000100000100001000100011101000011",
--  (468) multiplication_with_reduction_242
-- reg_a = o2_X; reg_b = prime7; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011101010111",
--  (469) multiplication_with_reduction_243
-- reg_a = a3_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011001100011",
--  (470) multiplication_with_reduction_244
-- reg_a = o3_X; reg_b = prime6; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011001110111",
--  (471) multiplication_with_reduction_245
-- reg_a = a4_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010110000011",
--  (472) multiplication_with_reduction_246
-- reg_a = o4_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010110010111",
--  (473) multiplication_with_reduction_247
-- reg_a = a5_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010010100011",
--  (474) multiplication_with_reduction_248
-- reg_a = o5_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010010110111",
--  (475) multiplication_with_reduction_249
-- reg_a = a6_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001111000011",
--  (476) multiplication_with_reduction_250
-- reg_a = o6_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001111010111",
--  (477) multiplication_with_reduction_251
-- reg_a = a7_X; reg_b = b2_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001111000000000100000000000100100001011100011",
--  (478) multiplication_with_reduction_252
-- reg_a = o7_X; reg_b = prime2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000001000101011110111",
--  (479) multiplication_with_reduction_253
-- reg_a = a3_X; reg_b = b7_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001111000000000100000100001000100011101100011",
--  (480) multiplication_with_reduction_254
-- reg_a = o3_X; reg_b = prime7; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011101110111",
--  (481) multiplication_with_reduction_255
-- reg_a = a4_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011010000011",
--  (482) multiplication_with_reduction_256
-- reg_a = o4_X; reg_b = prime6; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011010010111",
--  (483) multiplication_with_reduction_257
-- reg_a = a5_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010110100011",
--  (484) multiplication_with_reduction_258
-- reg_a = o5_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010110110111",
--  (485) multiplication_with_reduction_259
-- reg_a = a6_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010011000011",
--  (486) multiplication_with_reduction_260
-- reg_a = o6_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010011010111",
--  (487) multiplication_with_reduction_261
-- reg_a = a7_X; reg_b = b3_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001111000000000100000000000100100001111100011",
--  (488) multiplication_with_reduction_262
-- reg_a = o7_X; reg_b = prime3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000001101001111110111",
--  (489) multiplication_with_reduction_263
-- reg_a = a4_X; reg_b = b7_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001111000000000100000100001000100011110000011",
--  (490) multiplication_with_reduction_264
-- reg_a = o4_X; reg_b = prime7; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011110010111",
--  (491) multiplication_with_reduction_265
-- reg_a = a5_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011010100011",
--  (492) multiplication_with_reduction_266
-- reg_a = o5_X; reg_b = prime6; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011010110111",
--  (493) multiplication_with_reduction_267
-- reg_a = a6_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010111000011",
--  (494) multiplication_with_reduction_268
-- reg_a = o6_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010111010111",
--  (495) multiplication_with_reduction_269
-- reg_a = a7_X; reg_b = b4_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001111000000000100000000000100100010011100011",
--  (496) multiplication_with_reduction_270
-- reg_a = o7_X; reg_b = prime4; reg_acc = reg_o; o3_X = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000010001110011110111",
--  (497) multiplication_with_reduction_271
-- reg_a = a5_X; reg_b = b7_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001111000000000100000100001000100011110100011",
--  (498) multiplication_with_reduction_272
-- reg_a = o5_X; reg_b = prime7; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011110110111",
--  (499) multiplication_with_reduction_273
-- reg_a = a6_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011011000011",
--  (500) multiplication_with_reduction_274
-- reg_a = o6_X; reg_b = prime6; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011011010111",
--  (501) multiplication_with_reduction_275
-- reg_a = a7_X; reg_b = b5_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001111000000000100000000000100100010111100011",
--  (502) multiplication_with_reduction_276
-- reg_a = o7_X; reg_b = prime5; reg_acc = reg_o; o4_X = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000010110010111110111",
--  (503) multiplication_with_reduction_277
-- reg_a = a6_X; reg_b = b7_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001111000000000100000100001000100011111000011",
--  (504) multiplication_with_reduction_278
-- reg_a = o6_X; reg_b = prime7; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011111010111",
--  (505) multiplication_with_reduction_279
-- reg_a = a7_X; reg_b = b6_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001111000000000100000000000100100011011100011",
--  (506) multiplication_with_reduction_280
-- reg_a = o7_X; reg_b = prime6; reg_acc = reg_o; o5_X = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000011010111011110111",
--  (507) multiplication_with_reduction_281
-- reg_a = a7_X; reg_b = b7_X; reg_acc = reg_o >> 256; Enable sign a, b; operation : a*b + acc;
"000000100001111000000000100000100001100100011111100011",
--  (508) multiplication_with_reduction_282
-- reg_a = o7_X; reg_b = prime7; reg_acc = reg_o; o6_X = reg_o; o7_0 = reg_o >> 256; operation : a*b + acc;
"000000100001111001110000100000000000011111011111110111",
--  (509) multiplication_with_reduction_283
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (510) multiplication_with_reduction_special_prime_1_0
-- -- In case of size 1
-- reg_a = a0_X; reg_b = b0_X; reg_acc = 0; Enable sign a,b; operation : a*b + acc;
"000000100001000000000000100000010000000100000000000011",
--  (511) multiplication_with_reduction_special_prime_1_1
-- reg_a = 0; reg_b = 0; reg_acc = reg_o >> 256; o0_X = reg_o; operation : a*b + acc;
"000000100001000000010000100000101110000100000000000011",
--  (512) multiplication_with_reduction_special_prime_1_2
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (513) multiplication_with_reduction_special_prime_1_3
-- -- In case of sizes 2, 3, 4, 5, 6, 7, 8
-- reg_a = a0_X; reg_b = b0_X; reg_acc = 0; o0_X = reg_o; operation : a*b + acc;
"000011100001001000010000100000010000000100000000000011",
--  (514) multiplication_with_reduction_special_prime_1_4
-- -- In case of size 2
-- reg_a = a0_X; reg_b = b1_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001001000000000100000100001000100000100000011",
--  (515) multiplication_with_reduction_special_prime_1_5
-- reg_a = o0_X; reg_b = primeSP1; reg_acc = reg_o; operation : a*b + acc;
"000000100001001000000000100000000000000100000100010111",
--  (516) multiplication_with_reduction_special_prime_1_6
-- reg_a = a1_X; reg_b = b0_X; reg_acc = reg_o; o1_X = reg_o; Enable sign a; operation : a*b + acc;
"000000100001001000010000100000000000101000100000100011",
--  (517) multiplication_with_reduction_special_prime_1_7
-- reg_a = a1_X; reg_b = b1_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001001000000000100000100001100100000100100011",
--  (518) multiplication_with_reduction_special_prime_1_8
-- reg_a = o1_X; reg_b = primeSP1; reg_acc = reg_o; o0_X = reg_o; o1_X = reg_o >> 256; operation : a*b + acc;
"000000100001001001110000100000000000000100000100110111",
--  (519) multiplication_with_reduction_special_prime_1_9
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (520) multiplication_with_reduction_special_prime_1_10
-- -- In case of sizes 3, 4, 5, 6, 7, 8
-- reg_a = a0_X; reg_b = b1_X; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001010000000000100000100000000100000100000011",
--  (521) multiplication_with_reduction_special_prime_1_11
-- reg_a = o0_X; reg_b = primeSP1; reg_acc = reg_o; operation : a*b + acc;
"000000100001010000000000100000000000000100000100010111",
--  (522) multiplication_with_reduction_special_prime_1_12
-- reg_a = a1_X; reg_b = b0_X; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
"000000100001010000010000100000000000001000100000100011",
--  (523) multiplication_with_reduction_special_prime_1_13
-- reg_a = o0_X; reg_b = primeSP2; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001010000000000100000100000000100001000010111",
--  (524) multiplication_with_reduction_special_prime_1_14
-- reg_a = a1_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001010000000000100000000000000100000100100011",
--  (525) multiplication_with_reduction_special_prime_1_15
-- reg_a = o1_X; reg_b = primeSP1; reg_acc = reg_o; operation : a*b + acc;
"000101000001010000000000100000000000000100000100110111",
--  (526) multiplication_with_reduction_special_prime_1_16
-- -- In case of size 3
-- reg_a = a0_X; reg_b = b2_X; reg_acc = reg_o; Enable sign b; operation : a*b + acc;
"000000100001010000000000100000000001000100001000000011",
--  (527) multiplication_with_reduction_special_prime_1_17
-- reg_a = a2_X; reg_b = b0_X; reg_acc = reg_o; o2_X = reg_o; Enable sign a; operation : a*b + acc;
"000000100001010000010000100000000000101101000001000011",
--  (528) multiplication_with_reduction_special_prime_1_18
-- reg_a = a1_X; reg_b = b2_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001010000000000100000100001000100001000100011",
--  (529) multiplication_with_reduction_special_prime_1_19
-- reg_a = o1_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
"000000100001010000000000100000000000000100001000110111",
--  (530) multiplication_with_reduction_special_prime_1_20
-- reg_a = a2_X; reg_b = b1_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001010000000000100000000000100100000101000011",
--  (531) multiplication_with_reduction_special_prime_1_21
-- reg_a = o2_X; reg_b = primeSP1; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
"000000100001010000010000100000000000000100000101010111",
--  (532) multiplication_with_reduction_special_prime_1_22
-- reg_a = a2_X; reg_b = b2_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001010000000000100000100001100100001001000011",
--  (533) multiplication_with_reduction_special_prime_1_23
-- reg_a = o2_X; reg_b = primeSP2; reg_acc = reg_o; o1_X = reg_o; o2_X = reg_o >> 256; operation : a*b + acc;
"000000100001010001110000100000000000001000101001010111",
--  (534) multiplication_with_reduction_special_prime_1_24
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (535) multiplication_with_reduction_special_prime_1_25
-- -- In case of sizes 4, 5, 6, 7, 8
-- reg_a = a0_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001011000000000100000000000000100001000000011",
--  (536) multiplication_with_reduction_special_prime_1_26
-- reg_a = a2_X; reg_b = b0_X; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
"000000100001011000010000100000000000001101000001000011",
--  (537) multiplication_with_reduction_special_prime_1_27
-- reg_a = o0_X; reg_b = primeSP3; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001011000000000100000100000000100001100010111",
--  (538) multiplication_with_reduction_special_prime_1_28
-- reg_a = a1_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001011000000000100000000000000100001000100011",
--  (539) multiplication_with_reduction_special_prime_1_29
-- reg_a = o1_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
"000000100001011000000000100000000000000100001000110111",
--  (540) multiplication_with_reduction_special_prime_1_30
-- reg_a = a2_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001011000000000100000000000000100000101000011",
--  (541) multiplication_with_reduction_special_prime_1_31
-- reg_a = o2_X; reg_b = primeSP1; reg_acc = reg_o; operation : a*b + acc;
"001000000001011000000000100000000000000100000101010111",
--  (542) multiplication_with_reduction_special_prime_1_32
-- -- In case of size 4
-- reg_a = a0_X; reg_b = b3_X; reg_acc = reg_o; Enable sign b; operation : a*b + acc;
"000000100001011000000000100000000001000100001100000011",
--  (543) multiplication_with_reduction_special_prime_1_33
-- reg_a = a3_X; reg_b = b0_X; reg_acc = reg_o; o3_X = reg_o; Enable sign a; operation : a*b + acc;
"000000100001011000010000100000000000100001100001100011",
--  (544) multiplication_with_reduction_special_prime_1_34
-- reg_a = a1_X; reg_b = b3_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001011000000000100000100001000100001100100011",
--  (545) multiplication_with_reduction_special_prime_1_35
-- reg_a = o1_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001011000000000100000000000000100001100110111",
--  (546) multiplication_with_reduction_special_prime_1_36
-- reg_a = a2_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001011000000000100000000000000100001001000011",
--  (547) multiplication_with_reduction_special_prime_1_37
-- reg_a = o2_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
"000000100001011000000000100000000000000100001001010111",
--  (548) multiplication_with_reduction_special_prime_1_38
-- reg_a = a3_X; reg_b = b1_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001011000000000100000000000100100000101100011",
--  (549) multiplication_with_reduction_special_prime_1_39
-- reg_a = o3_X; reg_b = primeSP1; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
"000000100001011000010000100000000000000100000101110111",
--  (550) multiplication_with_reduction_special_prime_1_40
-- reg_a = a2_X; reg_b = b3_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001011000000000100000100001000100001101000011",
--  (551) multiplication_with_reduction_special_prime_1_41
-- reg_a = o2_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001011000000000100000000000000100001101010111",
--  (552) multiplication_with_reduction_special_prime_1_42
-- reg_a = a3_X; reg_b = b2_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001011000000000100000000000100100001001100011",
--  (553) multiplication_with_reduction_special_prime_1_43
-- reg_a = o3_X; reg_b = primeSP2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
"000000100001011000010000100000000000001000101001110111",
--  (554) multiplication_with_reduction_special_prime_1_44
-- reg_a = a3_X; reg_b = b3_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001011000000000100000100001100100001101100011",
--  (555) multiplication_with_reduction_special_prime_1_45
-- reg_a = o3_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; o3_X = reg_o >> 256; operation : a*b + acc;
"000000100001011001110000100000000000001101001101110111",
--  (556) multiplication_with_reduction_special_prime_1_46
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (557) multiplication_with_reduction_special_prime_1_47
-- -- In case of sizes 5, 6, 7, 8
-- reg_a = a0_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001100000011",
--  (558) multiplication_with_reduction_special_prime_1_48
-- reg_a = a3_X; reg_b = b0_X; reg_acc = reg_o; o3_X = reg_o; operation : a*b + acc;
"000000100001100000010000100000000000010001100001100011",
--  (559) multiplication_with_reduction_special_prime_1_49
-- reg_a = o0_X; reg_b = primeSP4; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001100000000000100000100000000100010000010111",
--  (560) multiplication_with_reduction_special_prime_1_50
-- reg_a = a1_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001100100011",
--  (561) multiplication_with_reduction_special_prime_1_51
-- reg_a = o1_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001100110111",
--  (562) multiplication_with_reduction_special_prime_1_52
-- reg_a = a2_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001001000011",
--  (563) multiplication_with_reduction_special_prime_1_53
-- reg_a = o2_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001001010111",
--  (564) multiplication_with_reduction_special_prime_1_54
-- reg_a = a3_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100000101100011",
--  (565) multiplication_with_reduction_special_prime_1_55
-- reg_a = o3_X; reg_b = primeSP1; reg_acc = reg_o; operation : a*b + acc;
"001100000001100000000000100000000000000100000101110111",
--  (566) multiplication_with_reduction_special_prime_1_56
-- -- In case of size 5
-- reg_a = a0_X; reg_b = b4_X; reg_acc = reg_o; Enable sign b; operation : a*b + acc;
"000000100001100000000000100000000001000100010000000011",
--  (567) multiplication_with_reduction_special_prime_1_57
-- reg_a = a4_X; reg_b = b0_X; reg_acc = reg_o; o4_X = reg_o; Enable sign a; operation : a*b + acc;
"000000100001100000010000100000000000110110000010000011",
--  (568) multiplication_with_reduction_special_prime_1_58
-- reg_a = a1_X; reg_b = b4_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001100000000000100000100001000100010000100011",
--  (569) multiplication_with_reduction_special_prime_1_59
-- reg_a = o1_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100010000110111",
--  (570) multiplication_with_reduction_special_prime_1_60
-- reg_a = a2_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001101000011",
--  (571) multiplication_with_reduction_special_prime_1_61
-- reg_a = o2_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001101010111",
--  (572) multiplication_with_reduction_special_prime_1_62
-- reg_a = a3_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001001100011",
--  (573) multiplication_with_reduction_special_prime_1_63
-- reg_a = o3_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001001110111",
--  (574) multiplication_with_reduction_special_prime_1_64
-- reg_a = a4_X; reg_b = b1_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001100000000000100000000000100100000110000011",
--  (575) multiplication_with_reduction_special_prime_1_65
-- reg_a = o4_X; reg_b = primeSP1; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
"000000100001100000010000100000000000000100000110010111",
--  (576) multiplication_with_reduction_special_prime_1_66
-- reg_a = a2_X; reg_b = b4_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001100000000000100000100001000100010001000011",
--  (577) multiplication_with_reduction_special_prime_1_67
-- reg_a = o2_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100010001010111",
--  (578) multiplication_with_reduction_special_prime_1_68
-- reg_a = a3_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001101100011",
--  (579) multiplication_with_reduction_special_prime_1_69
-- reg_a = o3_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001101110111",
--  (580) multiplication_with_reduction_special_prime_1_70
-- reg_a = a4_X; reg_b = b2_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001100000000000100000000000100100001010000011",
--  (581) multiplication_with_reduction_special_prime_1_71
-- reg_a = o4_X; reg_b = primeSP2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
"000000100001100000010000100000000000001000101010010111",
--  (582) multiplication_with_reduction_special_prime_1_72
-- reg_a = a3_X; reg_b = b4_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001100000000000100000100001000100010001100011",
--  (583) multiplication_with_reduction_special_prime_1_73
-- reg_a = o3_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100010001110111",
--  (584) multiplication_with_reduction_special_prime_1_74
-- reg_a = a4_X; reg_b = b3_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001100000000000100000000000100100001110000011",
--  (585) multiplication_with_reduction_special_prime_1_75
-- reg_a = o4_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
"000000100001100000010000100000000000001101001110010111",
--  (586) multiplication_with_reduction_special_prime_1_76
-- reg_a = a4_X; reg_b = b4_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001100000000000100000100001100100010010000011",
--  (587) multiplication_with_reduction_special_prime_1_77
-- reg_a = o4_X; reg_b = primeSP4; reg_acc = reg_o; o3_X = reg_o; o4_X = reg_o >> 256; operation : a*b + acc;
"000000100001100001110000100000000000010001110010010111",
--  (588) multiplication_with_reduction_special_prime_1_78
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (589) multiplication_with_reduction_special_prime_1_79
-- -- In case of sizes 6, 7, 8
-- reg_a = a0_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010000000011",
--  (590) multiplication_with_reduction_special_prime_1_80
-- reg_a = a4_X; reg_b = b0_X; reg_acc = reg_o; o4_X = reg_o; operation : a*b + acc;
"000000100001101000010000100000000000010110000010000011",
--  (591) multiplication_with_reduction_special_prime_1_81
-- reg_a = o0_X; reg_b = primeSP5; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001101000000000100000100000000100010100010111",
--  (592) multiplication_with_reduction_special_prime_1_82
-- reg_a = a1_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010000100011",
--  (593) multiplication_with_reduction_special_prime_1_83
-- reg_a = o1_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010000110111",
--  (594) multiplication_with_reduction_special_prime_1_84
-- reg_a = a2_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001101000011",
--  (595) multiplication_with_reduction_special_prime_1_85
-- reg_a = o2_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001101010111",
--  (596) multiplication_with_reduction_special_prime_1_86
-- reg_a = a3_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001001100011",
--  (597) multiplication_with_reduction_special_prime_1_87
-- reg_a = o3_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001001110111",
--  (598) multiplication_with_reduction_special_prime_1_88
-- reg_a = a4_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100000110000011",
--  (599) multiplication_with_reduction_special_prime_1_89
-- reg_a = o4_X; reg_b = primeSP1; reg_acc = reg_o; operation : a*b + acc;
"010001000001101000000000100000000000000100000110010111",
--  (600) multiplication_with_reduction_special_prime_1_90
-- -- In case of size 6
-- reg_a = a0_X; reg_b = b5_X; reg_acc = reg_o; Enable sign b; operation : a*b + acc;
"000000100001101000000000100000000001000100010100000011",
--  (601) multiplication_with_reduction_special_prime_1_91
-- reg_a = a5_X; reg_b = b0_X; reg_acc = reg_o; o5_X = reg_o; Enable sign a; operation : a*b + acc;
"000000100001101000010000100000000000111010100010100011",
--  (602) multiplication_with_reduction_special_prime_1_92
-- reg_a = a1_X; reg_b = b5_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001101000000000100000100001000100010100100011",
--  (603) multiplication_with_reduction_special_prime_1_93
-- reg_a = o1_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010100110111",
--  (604) multiplication_with_reduction_special_prime_1_94
-- reg_a = a2_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010001000011",
--  (605) multiplication_with_reduction_special_prime_1_95
-- reg_a = o2_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010001010111",
--  (606) multiplication_with_reduction_special_prime_1_96
-- reg_a = a3_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001101100011",
--  (607) multiplication_with_reduction_special_prime_1_97
-- reg_a = o3_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001101110111",
--  (608) multiplication_with_reduction_special_prime_1_98
-- reg_a = a4_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001010000011",
--  (609) multiplication_with_reduction_special_prime_1_99
-- reg_a = o4_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001010010111",
--  (610) multiplication_with_reduction_special_prime_1_100
-- reg_a = a5_X; reg_b = b1_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001101000000000100000000000100100000110100011",
--  (611) multiplication_with_reduction_special_prime_1_101
-- reg_a = o5_X; reg_b = primeSP1; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
"000000100001101000010000100000000000000100000110110111",
--  (612) multiplication_with_reduction_special_prime_1_102
-- reg_a = a2_X; reg_b = b5_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001101000000000100000100001000100010101000011",
--  (613) multiplication_with_reduction_special_prime_1_103
-- reg_a = o2_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010101010111",
--  (614) multiplication_with_reduction_special_prime_1_104
-- reg_a = a3_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010001100011",
--  (615) multiplication_with_reduction_special_prime_1_105
-- reg_a = o3_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010001110111",
--  (616) multiplication_with_reduction_special_prime_1_106
-- reg_a = a4_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001110000011",
--  (617) multiplication_with_reduction_special_prime_1_107
-- reg_a = o4_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001110010111",
--  (618) multiplication_with_reduction_special_prime_1_108
-- reg_a = a5_X; reg_b = b2_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001101000000000100000000000100100001010100011",
--  (619) multiplication_with_reduction_special_prime_1_109
-- reg_a = o5_X; reg_b = primeSP2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
"000000100001101000010000100000000000001000101010110111",
--  (620) multiplication_with_reduction_special_prime_1_110
-- reg_a = a3_X; reg_b = b5_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001101000000000100000100001000100010101100011",
--  (621) multiplication_with_reduction_special_prime_1_111
-- reg_a = o3_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010101110111",
--  (622) multiplication_with_reduction_special_prime_1_112
-- reg_a = a4_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010010000011",
--  (623) multiplication_with_reduction_special_prime_1_113
-- reg_a = o4_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010010010111",
--  (624) multiplication_with_reduction_special_prime_1_114
-- reg_a = a5_X; reg_b = b3_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001101000000000100000000000100100001110100011",
--  (625) multiplication_with_reduction_special_prime_1_115
-- reg_a = o5_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
"000000100001101000010000100000000000001101001110110111",
--  (626) multiplication_with_reduction_special_prime_1_116
-- reg_a = a4_X; reg_b = b5_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001101000000000100000100001000100010110000011",
--  (627) multiplication_with_reduction_special_prime_1_117
-- reg_a = o4_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010110010111",
--  (628) multiplication_with_reduction_special_prime_1_118
-- reg_a = a5_X; reg_b = b4_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001101000000000100000000000100100010010100011",
--  (629) multiplication_with_reduction_special_prime_1_119
-- reg_a = o5_X; reg_b = primeSP4; reg_acc = reg_o; o3_X = reg_o; operation : a*b + acc;
"000000100001101000010000100000000000010001110010110111",
--  (630) multiplication_with_reduction_special_prime_1_120
-- reg_a = a5_X; reg_b = b5_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001101000000000100000100001100100010110100011",
--  (631) multiplication_with_reduction_special_prime_1_121
-- reg_a = o5_X; reg_b = primeSP5; reg_acc = reg_o; o4_X = reg_o; o5_X = reg_o >> 256; operation : a*b + acc;
"000000100001101001110000100000000000010110010110110111",
--  (632) multiplication_with_reduction_special_prime_1_122
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (633) multiplication_with_reduction_special_prime_1_123
-- -- In case of sizes 7, 8
-- reg_a = a0_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010100000011",
--  (634) multiplication_with_reduction_special_prime_1_124
-- reg_a = a5_X; reg_b = b0_X; reg_acc = reg_o; o5_X = reg_o; operation : a*b + acc;
"000000100001110000010000100000000000011010100010100011",
--  (635) multiplication_with_reduction_special_prime_1_125
-- reg_a = o0_X; reg_b = primeSP6; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001110000000000100000100000000100011000010111",
--  (636) multiplication_with_reduction_special_prime_1_126
-- reg_a = a1_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010100100011",
--  (637) multiplication_with_reduction_special_prime_1_127
-- reg_a = o1_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010100110111",
--  (638) multiplication_with_reduction_special_prime_1_128
-- reg_a = a2_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010001000011",
--  (639) multiplication_with_reduction_special_prime_1_129
-- reg_a = o2_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010001010111",
--  (640) multiplication_with_reduction_special_prime_1_130
-- reg_a = a3_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001101100011",
--  (641) multiplication_with_reduction_special_prime_1_131
-- reg_a = o3_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001101110111",
--  (642) multiplication_with_reduction_special_prime_1_132
-- reg_a = a4_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001010000011",
--  (643) multiplication_with_reduction_special_prime_1_133
-- reg_a = o4_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001010010111",
--  (644) multiplication_with_reduction_special_prime_1_134
-- reg_a = a5_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100000110100011",
--  (645) multiplication_with_reduction_special_prime_1_135
-- reg_a = o5_X; reg_b = primeSP1; reg_acc = reg_o; operation : a*b + acc;
"010111000001110000000000100000000000000100000110110111",
--  (646) multiplication_with_reduction_special_prime_1_136
-- -- In case of size 7
-- reg_a = a0_X; reg_b = b6_X; reg_acc = reg_o; Enable sign b; operation : a*b + acc;
"000000100001110000000000100000000001000100011000000011",
--  (647) multiplication_with_reduction_special_prime_1_137
-- reg_a = a6_X; reg_b = b0_X; reg_acc = reg_o; o6_X = reg_o; Enable sign a; operation : a*b + acc;
"000000100001110000010000100000000000111111000011000011",
--  (648) multiplication_with_reduction_special_prime_1_138
-- reg_a = a1_X; reg_b = b6_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001110000000000100000100001000100011000100011",
--  (649) multiplication_with_reduction_special_prime_1_139
-- reg_a = o1_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100011000110111",
--  (650) multiplication_with_reduction_special_prime_1_140
-- reg_a = a2_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010101000011",
--  (651) multiplication_with_reduction_special_prime_1_141
-- reg_a = o2_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010101010111",
--  (652) multiplication_with_reduction_special_prime_1_142
-- reg_a = a3_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010001100011",
--  (653) multiplication_with_reduction_special_prime_1_143
-- reg_a = o3_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010001110111",
--  (654) multiplication_with_reduction_special_prime_1_144
-- reg_a = a4_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001110000011",
--  (655) multiplication_with_reduction_special_prime_1_145
-- reg_a = o4_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001110010111",
--  (656) multiplication_with_reduction_special_prime_1_146
-- reg_a = a5_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001010100011",
--  (657) multiplication_with_reduction_special_prime_1_147
-- reg_a = o5_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001010110111",
--  (658) multiplication_with_reduction_special_prime_1_148
-- reg_a = a6_X; reg_b = b1_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001110000000000100000000000100100000111000011",
--  (659) multiplication_with_reduction_special_prime_1_149
-- reg_a = o6_X; reg_b = primeSP1; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
"000000100001110000010000100000000000000100000111010111",
--  (660) multiplication_with_reduction_special_prime_1_150
-- reg_a = a2_X; reg_b = b6_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001110000000000100000100001000100011001000011",
--  (661) multiplication_with_reduction_special_prime_1_151
-- reg_a = o2_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100011001010111",
--  (662) multiplication_with_reduction_special_prime_1_152
-- reg_a = a3_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010101100011",
--  (663) multiplication_with_reduction_special_prime_1_153
-- reg_a = o3_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010101110111",
--  (664) multiplication_with_reduction_special_prime_1_154
-- reg_a = a4_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010010000011",
--  (665) multiplication_with_reduction_special_prime_1_155
-- reg_a = o4_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010010010111",
--  (666) multiplication_with_reduction_special_prime_1_156
-- reg_a = a5_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001110100011",
--  (667) multiplication_with_reduction_special_prime_1_157
-- reg_a = o5_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001110110111",
--  (668) multiplication_with_reduction_special_prime_1_158
-- reg_a = a6_X; reg_b = b2_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001110000000000100000000000100100001011000011",
--  (669) multiplication_with_reduction_special_prime_1_159
-- reg_a = o6_X; reg_b = primeSP2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
"000000100001110000010000100000000000001000101011010111",
--  (670) multiplication_with_reduction_special_prime_1_160
-- reg_a = a3_X; reg_b = b6_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001110000000000100000100001000100011001100011",
--  (671) multiplication_with_reduction_special_prime_1_161
-- reg_a = o3_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100011001110111",
--  (672) multiplication_with_reduction_special_prime_1_162
-- reg_a = a4_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010110000011",
--  (673) multiplication_with_reduction_special_prime_1_163
-- reg_a = o4_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010110010111",
--  (674) multiplication_with_reduction_special_prime_1_164
-- reg_a = a5_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010010100011",
--  (675) multiplication_with_reduction_special_prime_1_165
-- reg_a = o5_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010010110111",
--  (676) multiplication_with_reduction_special_prime_1_166
-- reg_a = a6_X; reg_b = b3_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001110000000000100000000000100100001111000011",
--  (677) multiplication_with_reduction_special_prime_1_167
-- reg_a = o6_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
"000000100001110000010000100000000000001101001111010111",
--  (678) multiplication_with_reduction_special_prime_1_168
-- reg_a = a4_X; reg_b = b6_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001110000000000100000100001000100011010000011",
--  (679) multiplication_with_reduction_special_prime_1_169
-- reg_a = o4_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100011010010111",
--  (680) multiplication_with_reduction_special_prime_1_170
-- reg_a = a5_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010110100011",
--  (681) multiplication_with_reduction_special_prime_1_171
-- reg_a = o5_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010110110111",
--  (682) multiplication_with_reduction_special_prime_1_172
-- reg_a = a6_X; reg_b = b4_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001110000000000100000000000100100010011000011",
--  (683) multiplication_with_reduction_special_prime_1_173
-- reg_a = o6_X; reg_b = primeSP4; reg_acc = reg_o; o3_X = reg_o; operation : a*b + acc;
"000000100001110000010000100000000000010001110011010111",
--  (684) multiplication_with_reduction_special_prime_1_174
-- reg_a = a5_X; reg_b = b6_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001110000000000100000100001000100011010100011",
--  (685) multiplication_with_reduction_special_prime_1_175
-- reg_a = o5_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100011010110111",
--  (686) multiplication_with_reduction_special_prime_1_176
-- reg_a = a6_X; reg_b = b5_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001110000000000100000000000100100010111000011",
--  (687) multiplication_with_reduction_special_prime_1_177
-- reg_a = o6_X; reg_b = primeSP5; reg_acc = reg_o; o4_X = reg_o; operation : a*b + acc;
"000000100001110000010000100000000000010110010111010111",
--  (688) multiplication_with_reduction_special_prime_1_178
-- reg_a = a6_X; reg_b = b6_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001110000000000100000100001100100011011000011",
--  (689) multiplication_with_reduction_special_prime_1_179
-- reg_a = o6_X; reg_b = primeSP6; reg_acc = reg_o; o5_X = reg_o; o6_X = reg_o >> 256; operation : a*b + acc;
"000000100001110001110000100000000000011010111011010111",
--  (690) multiplication_with_reduction_special_prime_1_180
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (691) multiplication_with_reduction_special_prime_1_181
-- -- In case of size 8
-- reg_a = a0_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011000000011",
--  (692) multiplication_with_reduction_special_prime_1_182
-- reg_a = a6_X; reg_b = b0_X; reg_acc = reg_o; o6_X = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000011111000011000011",
--  (693) multiplication_with_reduction_special_prime_1_183
-- reg_a = o0_X; reg_b = primeSP7; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001111000000000100000100000000100011100010111",
--  (694) multiplication_with_reduction_special_prime_1_184
-- reg_a = a1_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011000100011",
--  (695) multiplication_with_reduction_special_prime_1_185
-- reg_a = o1_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011000110111",
--  (696) multiplication_with_reduction_special_prime_1_186
-- reg_a = a2_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010101000011",
--  (697) multiplication_with_reduction_special_prime_1_187
-- reg_a = o2_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010101010111",
--  (698) multiplication_with_reduction_special_prime_1_188
-- reg_a = a3_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010001100011",
--  (699) multiplication_with_reduction_special_prime_1_189
-- reg_a = o3_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010001110111",
--  (700) multiplication_with_reduction_special_prime_1_190
-- reg_a = a4_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001110000011",
--  (701) multiplication_with_reduction_special_prime_1_191
-- reg_a = o4_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001110010111",
--  (702) multiplication_with_reduction_special_prime_1_192
-- reg_a = a5_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001010100011",
--  (703) multiplication_with_reduction_special_prime_1_193
-- reg_a = o5_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001010110111",
--  (704) multiplication_with_reduction_special_prime_1_194
-- reg_a = a6_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100000111000011",
--  (705) multiplication_with_reduction_special_prime_1_195
-- reg_a = o6_X; reg_b = primeSP1; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100000111010111",
--  (706) multiplication_with_reduction_special_prime_1_196
-- reg_a = a0_X; reg_b = b7_X; reg_acc = reg_o; Enable sign b; operation : a*b + acc;
"000000100001111000000000100000000001000100011100000011",
--  (707) multiplication_with_reduction_special_prime_1_197
-- reg_a = a7_X; reg_b = b0_X; reg_acc = reg_o; o7_X = reg_o; Enable sign a; operation : a*b + acc;
"000000100001111000010000100000000000100011100011100011",
--  (708) multiplication_with_reduction_special_prime_1_198
-- reg_a = a1_X; reg_b = b7_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001111000000000100000100001000100011100100011",
--  (709) multiplication_with_reduction_special_prime_1_199
-- reg_a = o1_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011100110111",
--  (710) multiplication_with_reduction_special_prime_1_200
-- reg_a = a2_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011001000011",
--  (711) multiplication_with_reduction_special_prime_1_201
-- reg_a = o2_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011001010111",
--  (712) multiplication_with_reduction_special_prime_1_202
-- reg_a = a3_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010101100011",
--  (713) multiplication_with_reduction_special_prime_1_203
-- reg_a = o3_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010101110111",
--  (714) multiplication_with_reduction_special_prime_1_204
-- reg_a = a4_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010010000011",
--  (715) multiplication_with_reduction_special_prime_1_205
-- reg_a = o4_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010010010111",
--  (716) multiplication_with_reduction_special_prime_1_206
-- reg_a = a5_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001110100011",
--  (717) multiplication_with_reduction_special_prime_1_207
-- reg_a = o5_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001110110111",
--  (718) multiplication_with_reduction_special_prime_1_208
-- reg_a = a6_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001011000011",
--  (719) multiplication_with_reduction_special_prime_1_209
-- reg_a = o6_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001011010111",
--  (720) multiplication_with_reduction_special_prime_1_210
-- reg_a = a7_X; reg_b = b1_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001111000000000100000000000100100000111100011",
--  (721) multiplication_with_reduction_special_prime_1_211
-- reg_a = o7_X; reg_b = primeSP1; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000000100000111110111",
--  (722) multiplication_with_reduction_special_prime_1_212
-- reg_a = a2_X; reg_b = b7_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001111000000000100000100001000100011101000011",
--  (723) multiplication_with_reduction_special_prime_1_213
-- reg_a = o2_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011101010111",
--  (724) multiplication_with_reduction_special_prime_1_214
-- reg_a = a3_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011001100011",
--  (725) multiplication_with_reduction_special_prime_1_215
-- reg_a = o3_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011001110111",
--  (726) multiplication_with_reduction_special_prime_1_216
-- reg_a = a4_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010110000011",
--  (727) multiplication_with_reduction_special_prime_1_217
-- reg_a = o4_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010110010111",
--  (728) multiplication_with_reduction_special_prime_1_218
-- reg_a = a5_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010010100011",
--  (729) multiplication_with_reduction_special_prime_1_219
-- reg_a = o5_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010010110111",
--  (730) multiplication_with_reduction_special_prime_1_220
-- reg_a = a6_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001111000011",
--  (731) multiplication_with_reduction_special_prime_1_221
-- reg_a = o6_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001111010111",
--  (732) multiplication_with_reduction_special_prime_1_222
-- reg_a = a7_X; reg_b = b2_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001111000000000100000000000100100001011100011",
--  (733) multiplication_with_reduction_special_prime_1_223
-- reg_a = o7_X; reg_b = primeSP2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000001000101011110111",
--  (734) multiplication_with_reduction_special_prime_1_224
-- reg_a = a3_X; reg_b = b7_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001111000000000100000100001000100011101100011",
--  (735) multiplication_with_reduction_special_prime_1_225
-- reg_a = o3_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011101110111",
--  (736) multiplication_with_reduction_special_prime_1_226
-- reg_a = a4_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011010000011",
--  (737) multiplication_with_reduction_special_prime_1_227
-- reg_a = o4_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011010010111",
--  (738) multiplication_with_reduction_special_prime_1_228
-- reg_a = a5_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010110100011",
--  (739) multiplication_with_reduction_special_prime_1_229
-- reg_a = o5_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010110110111",
--  (740) multiplication_with_reduction_special_prime_1_230
-- reg_a = a6_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010011000011",
--  (741) multiplication_with_reduction_special_prime_1_231
-- reg_a = o6_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010011010111",
--  (742) multiplication_with_reduction_special_prime_1_232
-- reg_a = a7_X; reg_b = b3_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001111000000000100000000000100100001111100011",
--  (743) multiplication_with_reduction_special_prime_1_233
-- reg_a = o7_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000001101001111110111",
--  (744) multiplication_with_reduction_special_prime_1_234
-- reg_a = a4_X; reg_b = b7_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001111000000000100000100001000100011110000011",
--  (745) multiplication_with_reduction_special_prime_1_235
-- reg_a = o4_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011110010111",
--  (746) multiplication_with_reduction_special_prime_1_236
-- reg_a = a5_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011010100011",
--  (747) multiplication_with_reduction_special_prime_1_237
-- reg_a = o5_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011010110111",
--  (748) multiplication_with_reduction_special_prime_1_238
-- reg_a = a6_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010111000011",
--  (749) multiplication_with_reduction_special_prime_1_239
-- reg_a = o6_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010111010111",
--  (750) multiplication_with_reduction_special_prime_1_240
-- reg_a = a7_X; reg_b = b4_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001111000000000100000000000100100010011100011",
--  (751) multiplication_with_reduction_special_prime_1_241
-- reg_a = o7_X; reg_b = primeSP4; reg_acc = reg_o; o3_X = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000010001110011110111",
--  (752) multiplication_with_reduction_special_prime_1_242
-- reg_a = a5_X; reg_b = b7_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001111000000000100000100001000100011110100011",
--  (753) multiplication_with_reduction_special_prime_1_243
-- reg_a = o5_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011110110111",
--  (754) multiplication_with_reduction_special_prime_1_244
-- reg_a = a6_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011011000011",
--  (755) multiplication_with_reduction_special_prime_1_245
-- reg_a = o6_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011011010111",
--  (756) multiplication_with_reduction_special_prime_1_246
-- reg_a = a7_X; reg_b = b5_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001111000000000100000000000100100010111100011",
--  (757) multiplication_with_reduction_special_prime_1_247
-- reg_a = o7_X; reg_b = primeSP5; reg_acc = reg_o; o4_X = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000010110010111110111",
--  (758) multiplication_with_reduction_special_prime_1_248
-- reg_a = a6_X; reg_b = b7_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001111000000000100000100001000100011111000011",
--  (759) multiplication_with_reduction_special_prime_1_249
-- reg_a = o6_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011111010111",
--  (760) multiplication_with_reduction_special_prime_1_250
-- reg_a = a7_X; reg_b = b6_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001111000000000100000000000100100011011100011",
--  (761) multiplication_with_reduction_special_prime_1_251
-- reg_a = o7_X; reg_b = primeSP6; reg_acc = reg_o; o5_X = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000011010111011110111",
--  (762) multiplication_with_reduction_special_prime_1_252
-- reg_a = a7_X; reg_b = b7_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001111000000000100000100001100100011111100011",
--  (763) multiplication_with_reduction_special_prime_1_253
-- reg_a = o7_X; reg_b = primeSP7; reg_acc = reg_o; o6_X = reg_o; o7_X = reg_o >> 256; operation : a*b + acc;
"000000100001111001110000100000000000011111011111110111",
--  (764) multiplication_with_reduction_special_prime_1_254
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (765) multiplication_with_reduction_special_prime_2_0
-- With 2 zeroes in prime sharp
-- -- In case of sizes 2, 3, 4, 5, 6, 7, 8
-- reg_a = a0_X; reg_b = b0_X; reg_acc = 0; o0_X = reg_o; operation : a*b + acc;
"000010100001001000010000100000010000000100000000000011",
--  (766) multiplication_with_reduction_special_prime_2_1
-- -- In case of size 2
-- reg_a = a0_X; reg_b = b1_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001001000000000100000100001000100000100000011",
--  (767) multiplication_with_reduction_special_prime_2_2
-- reg_a = a1_X; reg_b = b0_X; reg_acc = reg_o; o1_X = reg_o; Enable sign a; operation : a*b + acc;
"000000100001001000010000100000000000101000100000100011",
--  (768) multiplication_with_reduction_special_prime_2_3
-- reg_a = a1_X; reg_b = b1_X; reg_acc = reg_o >> 256; o0_X = reg_o; o1_X = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001001001110000100000100001100100000100100011",
--  (769) multiplication_with_reduction_special_prime_2_4
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (770) multiplication_with_reduction_special_prime_2_5
-- -- In case of sizes 3, 4, 5, 6, 7, 8
-- reg_a = a0_X; reg_b = b1_X; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001010000000000100000100000000100000100000011",
--  (771) multiplication_with_reduction_special_prime_2_6
-- reg_a = a1_X; reg_b = b0_X; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
"000000100001010000010000100000000000001000100000100011",
--  (772) multiplication_with_reduction_special_prime_2_7
-- reg_a = o0_X; reg_b = primeSP2; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001010000000000100000100000000100001000010111",
--  (773) multiplication_with_reduction_special_prime_2_8
-- reg_a = a1_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
"000100100001010000000000100000000000000100000100100011",
--  (774) multiplication_with_reduction_special_prime_2_9
-- -- In case of size 3
-- reg_a = a0_X; reg_b = b2_X; reg_acc = reg_o; Enable sign b; operation : a*b + acc;
"000000100001010000000000100000000001000100001000000011",
--  (775) multiplication_with_reduction_special_prime_2_10
-- reg_a = a2_X; reg_b = b0_X; reg_acc = reg_o; o2_X = reg_o; Enable sign a; operation : a*b + acc;
"000000100001010000010000100000000000101101000001000011",
--  (776) multiplication_with_reduction_special_prime_2_11
-- reg_a = a1_X; reg_b = b2_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001010000000000100000100001000100001000100011",
--  (777) multiplication_with_reduction_special_prime_2_12
-- reg_a = o1_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
"000000100001010000000000100000000000000100001000110111",
--  (778) multiplication_with_reduction_special_prime_2_13
-- reg_a = a2_X; reg_b = b1_X; reg_acc = reg_o; Enable sign a; o0_X = reg_o; operation : a*b + acc;
"000000100001010000010000100000000000100100000101000011",
--  (779) multiplication_with_reduction_special_prime_2_14
-- reg_a = a2_X; reg_b = b2_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001010000000000100000100001100100001001000011",
--  (780) multiplication_with_reduction_special_prime_2_15
-- reg_a = o2_X; reg_b = primeSP2; reg_acc = reg_o; o1_X = reg_o; o2_X = reg_o >> 256; operation : a*b + acc;
"000000100001010001110000100000000000001000101001010111",
--  (781) multiplication_with_reduction_special_prime_2_16
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (782) multiplication_with_reduction_special_prime_2_17
-- -- In case of sizes 4, 5, 6, 7, 8
-- reg_a = a0_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001011000000000100000000000000100001000000011",
--  (783) multiplication_with_reduction_special_prime_2_18
-- reg_a = a2_X; reg_b = b0_X; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
"000000100001011000010000100000000000001101000001000011",
--  (784) multiplication_with_reduction_special_prime_2_19
-- reg_a = o0_X; reg_b = primeSP3; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001011000000000100000100000000100001100010111",
--  (785) multiplication_with_reduction_special_prime_2_20
-- reg_a = a1_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001011000000000100000000000000100001000100011",
--  (786) multiplication_with_reduction_special_prime_2_21
-- reg_a = o1_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
"000000100001011000000000100000000000000100001000110111",
--  (787) multiplication_with_reduction_special_prime_2_22
-- reg_a = a2_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
"000111100001011000000000100000000000000100000101000011",
--  (788) multiplication_with_reduction_special_prime_2_23
-- -- In case of size 4
-- reg_a = a0_X; reg_b = b3_X; reg_acc = reg_o; Enable sign b; operation : a*b + acc;
"000000100001011000000000100000000001000100001100000011",
--  (789) multiplication_with_reduction_special_prime_2_24
-- reg_a = a3_X; reg_b = b0_X; reg_acc = reg_o; o3_X = reg_o; Enable sign a; operation : a*b + acc;
"000000100001011000010000100000000000100001100001100011",
--  (790) multiplication_with_reduction_special_prime_2_25
-- reg_a = a1_X; reg_b = b3_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001011000000000100000100001000100001100100011",
--  (791) multiplication_with_reduction_special_prime_2_26
-- reg_a = o1_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001011000000000100000000000000100001100110111",
--  (792) multiplication_with_reduction_special_prime_2_27
-- reg_a = a2_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001011000000000100000000000000100001001000011",
--  (793) multiplication_with_reduction_special_prime_2_28
-- reg_a = o2_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
"000000100001011000000000100000000000000100001001010111",
--  (794) multiplication_with_reduction_special_prime_2_29
-- reg_a = a3_X; reg_b = b1_X; reg_acc = reg_o; Enable sign a; o0_X = reg_o; operation : a*b + acc;
"000000100001011000010000100000000000100100000101100011",
--  (795) multiplication_with_reduction_special_prime_2_30
-- reg_a = a2_X; reg_b = b3_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001011000000000100000100001000100001101000011",
--  (796) multiplication_with_reduction_special_prime_2_31
-- reg_a = o2_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001011000000000100000000000000100001101010111",
--  (797) multiplication_with_reduction_special_prime_2_32
-- reg_a = a3_X; reg_b = b2_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001011000000000100000000000100100001001100011",
--  (798) multiplication_with_reduction_special_prime_2_33
-- reg_a = o3_X; reg_b = primeSP2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
"000000100001011000010000100000000000001000101001110111",
--  (799) multiplication_with_reduction_special_prime_2_34
-- reg_a = a3_X; reg_b = b3_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001011000000000100000100001100100001101100011",
--  (800) multiplication_with_reduction_special_prime_2_35
-- reg_a = o3_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; o3_X = reg_o >> 256; operation : a*b + acc;
"000000100001011001110000100000000000001101001101110111",
--  (801) multiplication_with_reduction_special_prime_2_36
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (802) multiplication_with_reduction_special_prime_2_37
-- -- In case of sizes 5, 6, 7, 8
-- reg_a = a0_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001100000011",
--  (803) multiplication_with_reduction_special_prime_2_38
-- reg_a = a3_X; reg_b = b0_X; reg_acc = reg_o; o3_X = reg_o; operation : a*b + acc;
"000000100001100000010000100000000000010001100001100011",
--  (804) multiplication_with_reduction_special_prime_2_39
-- reg_a = o0_X; reg_b = primeSP4; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001100000000000100000100000000100010000010111",
--  (805) multiplication_with_reduction_special_prime_2_40
-- reg_a = a1_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001100100011",
--  (806) multiplication_with_reduction_special_prime_2_41
-- reg_a = o1_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001100110111",
--  (807) multiplication_with_reduction_special_prime_2_42
-- reg_a = a2_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001001000011",
--  (808) multiplication_with_reduction_special_prime_2_43
-- reg_a = o2_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001001010111",
--  (809) multiplication_with_reduction_special_prime_2_44
-- reg_a = a3_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
"001011100001100000000000100000000000000100000101100011",
--  (810) multiplication_with_reduction_special_prime_2_45
-- In case of size 5
-- reg_a = a0_X; reg_b = b4_X; reg_acc = reg_o; Enable sign b; operation : a*b + acc;
"000000100001100000000000100000000001000100010000000011",
--  (811) multiplication_with_reduction_special_prime_2_46
-- reg_a = a4_X; reg_b = b0_X; reg_acc = reg_o; o4_X = reg_o; Enable sign a; operation : a*b + acc;
"000000100001100000010000100000000000100010000010000011",
--  (812) multiplication_with_reduction_special_prime_2_47
-- reg_a = a1_X; reg_b = b4_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001100000000000100000100001000100010000100011",
--  (813) multiplication_with_reduction_special_prime_2_48
-- reg_a = o1_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100010000110111",
--  (814) multiplication_with_reduction_special_prime_2_49
-- reg_a = a2_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001101000011",
--  (815) multiplication_with_reduction_special_prime_2_50
-- reg_a = o2_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001101010111",
--  (816) multiplication_with_reduction_special_prime_2_51
-- reg_a = a3_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001001100011",
--  (817) multiplication_with_reduction_special_prime_2_52
-- reg_a = o3_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001001110111",
--  (818) multiplication_with_reduction_special_prime_2_53
-- reg_a = a4_X; reg_b = b1_X; reg_acc = reg_o; o0_X = reg_o; Enable sign a; operation : a*b + acc;
"000000100001100000010000100000000000100100000110000011",
--  (819) multiplication_with_reduction_special_prime_2_54
-- reg_a = a2_X; reg_b = b4_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001100000000000100000100001000100010001000011",
--  (820) multiplication_with_reduction_special_prime_2_55
-- reg_a = o2_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100010001010111",
--  (821) multiplication_with_reduction_special_prime_2_56
-- reg_a = a3_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001101100011",
--  (822) multiplication_with_reduction_special_prime_2_57
-- reg_a = o3_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001101110111",
--  (823) multiplication_with_reduction_special_prime_2_58
-- reg_a = a4_X; reg_b = b2_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001100000000000100000000000100100001010000011",
--  (824) multiplication_with_reduction_special_prime_2_59
-- reg_a = o4_X; reg_b = primeSP2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
"000000100001100000010000100000000000001000101010010111",
--  (825) multiplication_with_reduction_special_prime_2_60
-- reg_a = a3_X; reg_b = b4_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001100000000000100000100001000100010001100011",
--  (826) multiplication_with_reduction_special_prime_2_61
-- reg_a = o3_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100010001110111",
--  (827) multiplication_with_reduction_special_prime_2_62
-- reg_a = a4_X; reg_b = b3_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001100000000000100000000000100100001110000011",
--  (828) multiplication_with_reduction_special_prime_2_63
-- reg_a = o4_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
"000000100001100000010000100000000000001101001110010111",
--  (829) multiplication_with_reduction_special_prime_2_64
-- reg_a = a4_X; reg_b = b4_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001100000000000100000100001100100010010000011",
--  (830) multiplication_with_reduction_special_prime_2_65
-- reg_a = o4_X; reg_b = primeSP4; reg_acc = reg_o; o3_X = reg_o; o4_X = reg_o >> 256; operation : a*b + acc;
"000000100001100001110000100000000000010001110010010111",
--  (831) multiplication_with_reduction_special_prime_2_66
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (832) multiplication_with_reduction_special_prime_2_67
-- -- In case of sizes 6, 7, 8
-- reg_a = a0_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010000000011",
--  (833) multiplication_with_reduction_special_prime_2_68
-- reg_a = a4_X; reg_b = b0_X; reg_acc = reg_o; o4_X = reg_o; operation : a*b + acc;
"000000100001101000010000100000000000010010000010000011",
--  (834) multiplication_with_reduction_special_prime_2_69
-- reg_a = o0_X; reg_b = primeSP5; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001101000000000100000100000000100010100010111",
--  (835) multiplication_with_reduction_special_prime_2_70
-- reg_a = a1_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010000100011",
--  (836) multiplication_with_reduction_special_prime_2_71
-- reg_a = o1_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010000110111",
--  (837) multiplication_with_reduction_special_prime_2_72
-- reg_a = a2_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001101000011",
--  (838) multiplication_with_reduction_special_prime_2_73
-- reg_a = o2_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001101010111",
--  (839) multiplication_with_reduction_special_prime_2_74
-- reg_a = a3_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001001100011",
--  (840) multiplication_with_reduction_special_prime_2_75
-- reg_a = o3_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001001110111",
--  (841) multiplication_with_reduction_special_prime_2_76
-- reg_a = a4_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
"010000100001101000000000100000000000000100000110000011",
--  (842) multiplication_with_reduction_special_prime_2_77
-- In case of size 6
-- reg_a = a0_X; reg_b = b5_X; reg_acc = reg_o; Enable sign b; operation : a*b + acc;
"000000100001101000000000100000000001000100010100000011",
--  (843) multiplication_with_reduction_special_prime_2_78
-- reg_a = a5_X; reg_b = b0_X; reg_acc = reg_o; o5_X = reg_o; Enable sign a; operation : a*b + acc;
"000000100001101000010000100000000000100010100010100011",
--  (844) multiplication_with_reduction_special_prime_2_79
-- reg_a = a1_X; reg_b = b5_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001101000000000100000100001000100010100100011",
--  (845) multiplication_with_reduction_special_prime_2_80
-- reg_a = o1_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010100110111",
--  (846) multiplication_with_reduction_special_prime_2_81
-- reg_a = a2_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010001000011",
--  (847) multiplication_with_reduction_special_prime_2_82
-- reg_a = o2_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010001010111",
--  (848) multiplication_with_reduction_special_prime_2_83
-- reg_a = a3_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001101100011",
--  (849) multiplication_with_reduction_special_prime_2_84
-- reg_a = o3_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001101110111",
--  (850) multiplication_with_reduction_special_prime_2_85
-- reg_a = a4_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001010000011",
--  (851) multiplication_with_reduction_special_prime_2_86
-- reg_a = o4_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001010010111",
--  (852) multiplication_with_reduction_special_prime_2_87
-- reg_a = a5_X; reg_b = b1_X; reg_acc = reg_o; o0_X = reg_o; Enable sign a; operation : a*b + acc;
"000000100001101000010000100000000000100100000110100011",
--  (853) multiplication_with_reduction_special_prime_2_88
-- reg_a = a2_X; reg_b = b5_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001101000000000100000100001000100010101000011",
--  (854) multiplication_with_reduction_special_prime_2_89
-- reg_a = o2_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010101010111",
--  (855) multiplication_with_reduction_special_prime_2_90
-- reg_a = a3_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010001100011",
--  (856) multiplication_with_reduction_special_prime_2_91
-- reg_a = o3_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010001110111",
--  (857) multiplication_with_reduction_special_prime_2_92
-- reg_a = a4_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001110000011",
--  (858) multiplication_with_reduction_special_prime_2_93
-- reg_a = o4_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001110010111",
--  (859) multiplication_with_reduction_special_prime_2_94
-- reg_a = a5_X; reg_b = b2_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001101000000000100000000000100100001010100011",
--  (860) multiplication_with_reduction_special_prime_2_95
-- reg_a = o5_X; reg_b = primeSP2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
"000000100001101000010000100000000000001000101010110111",
--  (861) multiplication_with_reduction_special_prime_2_96
-- reg_a = a3_X; reg_b = b5_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001101000000000100000100001000100010101100011",
--  (862) multiplication_with_reduction_special_prime_2_97
-- reg_a = o3_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010101110111",
--  (863) multiplication_with_reduction_special_prime_2_98
-- reg_a = a4_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010010000011",
--  (864) multiplication_with_reduction_special_prime_2_99
-- reg_a = o4_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010010010111",
--  (865) multiplication_with_reduction_special_prime_2_100
-- reg_a = a5_X; reg_b = b3_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001101000000000100000000000100100001110100011",
--  (866) multiplication_with_reduction_special_prime_2_101
-- reg_a = o5_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
"000000100001101000010000100000000000001101001110110111",
--  (867) multiplication_with_reduction_special_prime_2_102
-- reg_a = a4_X; reg_b = b5_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001101000000000100000100001000100010110000011",
--  (868) multiplication_with_reduction_special_prime_2_103
-- reg_a = o4_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010110010111",
--  (869) multiplication_with_reduction_special_prime_2_104
-- reg_a = a5_X; reg_b = b4_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001101000000000100000000000100100010010100011",
--  (870) multiplication_with_reduction_special_prime_2_105
-- reg_a = o5_X; reg_b = primeSP4; reg_acc = reg_o; o3_X = reg_o; operation : a*b + acc;
"000000100001101000010000100000000000010001110010110111",
--  (871) multiplication_with_reduction_special_prime_2_106
-- reg_a = a5_X; reg_b = b5_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001101000000000100000100001100100010110100011",
--  (872) multiplication_with_reduction_special_prime_2_107
-- reg_a = o5_X; reg_b = primeSP5; reg_acc = reg_o; o4_X = reg_o; o5_X = reg_o >> 256; operation : a*b + acc;
"000000100001101001110000100000000000010110010110110111",
--  (873) multiplication_with_reduction_special_prime_2_108
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (874) multiplication_with_reduction_special_prime_2_109
-- -- In case of sizes 7, 8
-- reg_a = a0_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010100000011",
--  (875) multiplication_with_reduction_special_prime_2_110
-- reg_a = a5_X; reg_b = b0_X; reg_acc = reg_o; o5_X = reg_o; operation : a*b + acc;
"000000100001110000010000100000000000011010100010100011",
--  (876) multiplication_with_reduction_special_prime_2_111
-- reg_a = o0_X; reg_b = primeSP6; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001110000000000100000100000000100011000010111",
--  (877) multiplication_with_reduction_special_prime_2_112
-- reg_a = a1_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010100100011",
--  (878) multiplication_with_reduction_special_prime_2_113
-- reg_a = o1_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010100110111",
--  (879) multiplication_with_reduction_special_prime_2_114
-- reg_a = a2_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010001000011",
--  (880) multiplication_with_reduction_special_prime_2_115
-- reg_a = o2_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010001010111",
--  (881) multiplication_with_reduction_special_prime_2_116
-- reg_a = a3_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001101100011",
--  (882) multiplication_with_reduction_special_prime_2_117
-- reg_a = o3_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001101110111",
--  (883) multiplication_with_reduction_special_prime_2_118
-- reg_a = a4_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001010000011",
--  (884) multiplication_with_reduction_special_prime_2_119
-- reg_a = o4_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001010010111",
--  (885) multiplication_with_reduction_special_prime_2_120
-- reg_a = a5_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
"010110100001110000000000100000000000000100000110100011",
--  (886) multiplication_with_reduction_special_prime_2_121
-- -- In case of size 7
-- reg_a = a0_X; reg_b = b6_X; reg_acc = reg_o; Enable sign b; operation : a*b + acc;
"000000100001110000000000100000000001000100011000000011",
--  (887) multiplication_with_reduction_special_prime_2_122
-- reg_a = a6_X; reg_b = b0_X; reg_acc = reg_o; o6_X = reg_o; Enable sign a; operation : a*b + acc;
"000000100001110000010000100000000000100011000011000011",
--  (888) multiplication_with_reduction_special_prime_2_123
-- reg_a = a1_X; reg_b = b6_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001110000000000100000100001000100011000100011",
--  (889) multiplication_with_reduction_special_prime_2_124
-- reg_a = o1_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100011000110111",
--  (890) multiplication_with_reduction_special_prime_2_125
-- reg_a = a2_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010101000011",
--  (891) multiplication_with_reduction_special_prime_2_126
-- reg_a = o2_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010101010111",
--  (892) multiplication_with_reduction_special_prime_2_127
-- reg_a = a3_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010001100011",
--  (893) multiplication_with_reduction_special_prime_2_128
-- reg_a = o3_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010001110111",
--  (894) multiplication_with_reduction_special_prime_2_129
-- reg_a = a4_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001110000011",
--  (895) multiplication_with_reduction_special_prime_2_130
-- reg_a = o4_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001110010111",
--  (896) multiplication_with_reduction_special_prime_2_131
-- reg_a = a5_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001010100011",
--  (897) multiplication_with_reduction_special_prime_2_132
-- reg_a = o5_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001010110111",
--  (898) multiplication_with_reduction_special_prime_2_133
-- reg_a = a6_X; reg_b = b1_X; reg_acc = reg_o; Enable sign a; o0_X = reg_o; operation : a*b + acc;
"000000100001110000010000100000000000100100000111000011",
--  (899) multiplication_with_reduction_special_prime_2_134
-- reg_a = a2_X; reg_b = b6_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001110000000000100000100001000100011001000011",
--  (900) multiplication_with_reduction_special_prime_2_135
-- reg_a = o2_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100011001010111",
--  (901) multiplication_with_reduction_special_prime_2_136
-- reg_a = a3_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010101100011",
--  (902) multiplication_with_reduction_special_prime_2_137
-- reg_a = o3_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010101110111",
--  (903) multiplication_with_reduction_special_prime_2_138
-- reg_a = a4_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010010000011",
--  (904) multiplication_with_reduction_special_prime_2_139
-- reg_a = o4_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010010010111",
--  (905) multiplication_with_reduction_special_prime_2_140
-- reg_a = a5_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001110100011",
--  (906) multiplication_with_reduction_special_prime_2_141
-- reg_a = o5_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001110110111",
--  (907) multiplication_with_reduction_special_prime_2_142
-- reg_a = a6_X; reg_b = b2_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001110000000000100000000000100100001011000011",
--  (908) multiplication_with_reduction_special_prime_2_143
-- reg_a = o6_X; reg_b = primeSP2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
"000000100001110000010000100000000000001000101011010111",
--  (909) multiplication_with_reduction_special_prime_2_144
-- reg_a = a3_X; reg_b = b6_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001110000000000100000100001000100011001100011",
--  (910) multiplication_with_reduction_special_prime_2_145
-- reg_a = o3_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100011001110111",
--  (911) multiplication_with_reduction_special_prime_2_146
-- reg_a = a4_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010110000011",
--  (912) multiplication_with_reduction_special_prime_2_147
-- reg_a = o4_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010110010111",
--  (913) multiplication_with_reduction_special_prime_2_148
-- reg_a = a5_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010010100011",
--  (914) multiplication_with_reduction_special_prime_2_149
-- reg_a = o5_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010010110111",
--  (915) multiplication_with_reduction_special_prime_2_150
-- reg_a = a6_X; reg_b = b3_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001110000000000100000000000100100001111000011",
--  (916) multiplication_with_reduction_special_prime_2_151
-- reg_a = o6_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
"000000100001110000010000100000000000001101001111010111",
--  (917) multiplication_with_reduction_special_prime_2_152
-- reg_a = a4_X; reg_b = b6_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001110000000000100000100001000100011010000011",
--  (918) multiplication_with_reduction_special_prime_2_153
-- reg_a = o4_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100011010010111",
--  (919) multiplication_with_reduction_special_prime_2_154
-- reg_a = a5_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010110100011",
--  (920) multiplication_with_reduction_special_prime_2_155
-- reg_a = o5_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010110110111",
--  (921) multiplication_with_reduction_special_prime_2_156
-- reg_a = a6_X; reg_b = b4_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001110000000000100000000000100100010011000011",
--  (922) multiplication_with_reduction_special_prime_2_157
-- reg_a = o6_X; reg_b = primeSP4; reg_acc = reg_o; o3_X = reg_o; operation : a*b + acc;
"000000100001110000010000100000000000010001110011010111",
--  (923) multiplication_with_reduction_special_prime_2_158
-- reg_a = a5_X; reg_b = b6_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001110000000000100000100001000100011010100011",
--  (924) multiplication_with_reduction_special_prime_2_159
-- reg_a = o5_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100011010110111",
--  (925) multiplication_with_reduction_special_prime_2_160
-- reg_a = a6_X; reg_b = b5_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001110000000000100000000000100100010111000011",
--  (926) multiplication_with_reduction_special_prime_2_161
-- reg_a = o6_X; reg_b = primeSP5; reg_acc = reg_o; o4_X = reg_o; operation : a*b + acc;
"000000100001110000010000100000000000010110010111010111",
--  (927) multiplication_with_reduction_special_prime_2_162
-- reg_a = a6_X; reg_b = b6_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001110000000000100000100001100100011011000011",
--  (928) multiplication_with_reduction_special_prime_2_163
-- reg_a = o6_X; reg_b = primeSP6; reg_acc = reg_o; o5_X = reg_o; o6_X = reg_o >> 256; operation : a*b + acc;
"000000100001110001110000100000000000011010111011010111",
--  (929) multiplication_with_reduction_special_prime_2_164
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (930) multiplication_with_reduction_special_prime_2_165
-- -- In case of size 8
-- reg_a = a0_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011000000011",
--  (931) multiplication_with_reduction_special_prime_2_166
-- reg_a = a6_X; reg_b = b0_X; reg_acc = reg_o; o6_X = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000011011000011000011",
--  (932) multiplication_with_reduction_special_prime_2_167
-- reg_a = o0_X; reg_b = primeSP7; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001111000000000100000100000000100011100010111",
--  (933) multiplication_with_reduction_special_prime_2_168
-- reg_a = a1_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011000100011",
--  (934) multiplication_with_reduction_special_prime_2_169
-- reg_a = o1_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011000110111",
--  (935) multiplication_with_reduction_special_prime_2_170
-- reg_a = a2_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010101000011",
--  (936) multiplication_with_reduction_special_prime_2_171
-- reg_a = o2_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010101010111",
--  (937) multiplication_with_reduction_special_prime_2_172
-- reg_a = a3_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010001100011",
--  (938) multiplication_with_reduction_special_prime_2_173
-- reg_a = o3_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010001110111",
--  (939) multiplication_with_reduction_special_prime_2_174
-- reg_a = a4_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001110000011",
--  (940) multiplication_with_reduction_special_prime_2_175
-- reg_a = o4_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001110010111",
--  (941) multiplication_with_reduction_special_prime_2_176
-- reg_a = a5_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001010100011",
--  (942) multiplication_with_reduction_special_prime_2_177
-- reg_a = o5_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001010110111",
--  (943) multiplication_with_reduction_special_prime_2_178
-- reg_a = a6_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100000111000011",
--  (944) multiplication_with_reduction_special_prime_2_179
-- reg_a = a0_X; reg_b = b7_X; reg_acc = reg_o; Enable sign b; operation : a*b + acc;
"000000100001111000000000100000000001000100011100000011",
--  (945) multiplication_with_reduction_special_prime_2_180
-- reg_a = a7_X; reg_b = b0_X; reg_acc = reg_o; o7_X = reg_o; Enable sign a; operation : a*b + acc;
"000000100001111000010000100000000000100011100011100011",
--  (946) multiplication_with_reduction_special_prime_2_181
-- reg_a = a1_X; reg_b = b7_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001111000000000100000100001000100011100100011",
--  (947) multiplication_with_reduction_special_prime_2_182
-- reg_a = o1_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011100110111",
--  (948) multiplication_with_reduction_special_prime_2_183
-- reg_a = a2_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011001000011",
--  (949) multiplication_with_reduction_special_prime_2_184
-- reg_a = o2_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011001010111",
--  (950) multiplication_with_reduction_special_prime_2_185
-- reg_a = a3_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010101100011",
--  (951) multiplication_with_reduction_special_prime_2_186
-- reg_a = o3_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010101110111",
--  (952) multiplication_with_reduction_special_prime_2_187
-- reg_a = a4_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010010000011",
--  (953) multiplication_with_reduction_special_prime_2_188
-- reg_a = o4_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010010010111",
--  (954) multiplication_with_reduction_special_prime_2_189
-- reg_a = a5_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001110100011",
--  (955) multiplication_with_reduction_special_prime_2_190
-- reg_a = o5_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001110110111",
--  (956) multiplication_with_reduction_special_prime_2_191
-- reg_a = a6_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001011000011",
--  (957) multiplication_with_reduction_special_prime_2_192
-- reg_a = o6_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001011010111",
--  (958) multiplication_with_reduction_special_prime_2_193
-- reg_a = a7_X; reg_b = b1_X; reg_acc = reg_o; Enable sign a; o0_X = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000100100000111100011",
--  (959) multiplication_with_reduction_special_prime_2_194
-- reg_a = a2_X; reg_b = b7_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001111000000000100000100001000100011101000011",
--  (960) multiplication_with_reduction_special_prime_2_195
-- reg_a = o2_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011101010111",
--  (961) multiplication_with_reduction_special_prime_2_196
-- reg_a = a3_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011001100011",
--  (962) multiplication_with_reduction_special_prime_2_197
-- reg_a = o3_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011001110111",
--  (963) multiplication_with_reduction_special_prime_2_198
-- reg_a = a4_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010110000011",
--  (964) multiplication_with_reduction_special_prime_2_199
-- reg_a = o4_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010110010111",
--  (965) multiplication_with_reduction_special_prime_2_200
-- reg_a = a5_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010010100011",
--  (966) multiplication_with_reduction_special_prime_2_201
-- reg_a = o5_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010010110111",
--  (967) multiplication_with_reduction_special_prime_2_202
-- reg_a = a6_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001111000011",
--  (968) multiplication_with_reduction_special_prime_2_203
-- reg_a = o6_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001111010111",
--  (969) multiplication_with_reduction_special_prime_2_204
-- reg_a = a7_X; reg_b = b2_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001111000000000100000000000100100001011100011",
--  (970) multiplication_with_reduction_special_prime_2_205
-- reg_a = o7_X; reg_b = primeSP2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000001000101011110111",
--  (971) multiplication_with_reduction_special_prime_2_206
-- reg_a = a3_X; reg_b = b7_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001111000000000100000100001000100011101100011",
--  (972) multiplication_with_reduction_special_prime_2_207
-- reg_a = o3_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011101110111",
--  (973) multiplication_with_reduction_special_prime_2_208
-- reg_a = a4_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011010000011",
--  (974) multiplication_with_reduction_special_prime_2_209
-- reg_a = o4_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011010010111",
--  (975) multiplication_with_reduction_special_prime_2_210
-- reg_a = a5_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010110100011",
--  (976) multiplication_with_reduction_special_prime_2_211
-- reg_a = o5_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010110110111",
--  (977) multiplication_with_reduction_special_prime_2_212
-- reg_a = a6_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010011000011",
--  (978) multiplication_with_reduction_special_prime_2_213
-- reg_a = o6_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010011010111",
--  (979) multiplication_with_reduction_special_prime_2_214
-- reg_a = a7_X; reg_b = b3_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001111000000000100000000000100100001111100011",
--  (980) multiplication_with_reduction_special_prime_2_215
-- reg_a = o7_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000001101001111110111",
--  (981) multiplication_with_reduction_special_prime_2_216
-- reg_a = a4_X; reg_b = b7_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001111000000000100000100001000100011110000011",
--  (982) multiplication_with_reduction_special_prime_2_217
-- reg_a = o4_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011110010111",
--  (983) multiplication_with_reduction_special_prime_2_218
-- reg_a = a5_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011010100011",
--  (984) multiplication_with_reduction_special_prime_2_219
-- reg_a = o5_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011010110111",
--  (985) multiplication_with_reduction_special_prime_2_220
-- reg_a = a6_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010111000011",
--  (986) multiplication_with_reduction_special_prime_2_221
-- reg_a = o6_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010111010111",
--  (987) multiplication_with_reduction_special_prime_2_222
-- reg_a = a7_X; reg_b = b4_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001111000000000100000000000100100010011100011",
--  (988) multiplication_with_reduction_special_prime_2_223
-- reg_a = o7_X; reg_b = primeSP4; reg_acc = reg_o; o3_X = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000010001110011110111",
--  (989) multiplication_with_reduction_special_prime_2_224
-- reg_a = a5_X; reg_b = b7_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001111000000000100000100001000100011110100011",
--  (990) multiplication_with_reduction_special_prime_2_225
-- reg_a = o5_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011110110111",
--  (991) multiplication_with_reduction_special_prime_2_226
-- reg_a = a6_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011011000011",
--  (992) multiplication_with_reduction_special_prime_2_227
-- reg_a = o6_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011011010111",
--  (993) multiplication_with_reduction_special_prime_2_228
-- reg_a = a7_X; reg_b = b5_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001111000000000100000000000100100010111100011",
--  (994) multiplication_with_reduction_special_prime_2_229
-- reg_a = o7_X; reg_b = primeSP5; reg_acc = reg_o; o4_X = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000010110010111110111",
--  (995) multiplication_with_reduction_special_prime_2_230
-- reg_a = a6_X; reg_b = b7_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001111000000000100000100001000100011111000011",
--  (996) multiplication_with_reduction_special_prime_2_231
-- reg_a = o6_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011111010111",
--  (997) multiplication_with_reduction_special_prime_2_232
-- reg_a = a7_X; reg_b = b6_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001111000000000100000000000100100011011100011",
--  (998) multiplication_with_reduction_special_prime_2_233
-- reg_a = o7_X; reg_b = primeSP6; reg_acc = reg_o; o5_X = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000011010111011110111",
--  (999) multiplication_with_reduction_special_prime_2_234
-- reg_a = a7_X; reg_b = b7_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001111000000000100000100001100100011111100011",
--  (1000) multiplication_with_reduction_special_prime_2_235
-- reg_a = o7_X; reg_b = primeSP7; reg_acc = reg_o; o6_X = reg_o; o7_X = reg_o >> 256; operation : a*b + acc;
"000000100001111001110000100000000000011111011111110111",
--  (1001) multiplication_with_reduction_special_prime_2_236
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (1002) multiplication_with_reduction_special_prime_3_0
-- -- In case of sizes 3, 4, 5, 6, 7, 8
-- reg_a = a0_X; reg_b = b0_X; reg_acc = 0; o0_X = reg_o; operation : a*b + acc;
"000000100001010000010000100000010000000100000000000011",
--  (1003) multiplication_with_reduction_special_prime_3_1
-- reg_a = a0_X; reg_b = b1_X; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001010000000000100000100000000100000100000011",
--  (1004) multiplication_with_reduction_special_prime_3_2
-- reg_a = a1_X; reg_b = b0_X; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
"000000100001010000010000100000000000001000100000100011",
--  (1005) multiplication_with_reduction_special_prime_3_3
-- reg_a = a1_X; reg_b = b1_X; reg_acc = reg_o >> 256; operation : a*b + acc;
"000011100001010000000000100000100000000100000100100011",
--  (1006) multiplication_with_reduction_special_prime_3_4
-- -- In case of size 3
-- reg_a = a0_X; reg_b = b2_X; reg_acc = reg_o; Enable sign b; operation : a*b + acc;
"000000100001010000000000100000000001000100001000000011",
--  (1007) multiplication_with_reduction_special_prime_3_5
-- reg_a = a2_X; reg_b = b0_X; reg_acc = reg_o; o2_X = reg_o; Enable sign a; operation : a*b + acc;
"000000100001010000010000100000000000101101000001000011",
--  (1008) multiplication_with_reduction_special_prime_3_6
-- reg_a = a1_X; reg_b = b2_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001010000000000100000100001000100001000100011",
--  (1009) multiplication_with_reduction_special_prime_3_7
-- reg_a = a2_X; reg_b = b1_X; reg_acc = reg_o; Enable sign a; o0_X = reg_o; operation : a*b + acc;
"000000100001010000010000100000000000100100000101000011",
--  (1010) multiplication_with_reduction_special_prime_3_8
-- reg_a = a2_X; reg_b = b2_X; reg_acc = reg_o >> 256; Enable sign a,b; o1_X = reg_o; o2_X = reg_o >> 256; operation : a*b + acc;
"000000100001010001110000100000100001100100001001000011",
--  (1011) multiplication_with_reduction_special_prime_3_9
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (1012) multiplication_with_reduction_special_prime_3_10
-- -- In case of sizes 4, 5, 6, 7, 8
-- reg_a = a0_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001011000000000100000000000000100001000000011",
--  (1013) multiplication_with_reduction_special_prime_3_11
-- reg_a = a2_X; reg_b = b0_X; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
"000000100001011000010000100000000000001101000001000011",
--  (1014) multiplication_with_reduction_special_prime_3_12
-- reg_a = o0_X; reg_b = primeSP3; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001011000000000100000100000000100001100010111",
--  (1015) multiplication_with_reduction_special_prime_3_13
-- reg_a = a1_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001011000000000100000000000000100001000100011",
--  (1016) multiplication_with_reduction_special_prime_3_14
-- reg_a = a2_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
"000110100001011000000000100000000000000100000101000011",
--  (1017) multiplication_with_reduction_special_prime_3_15
-- -- In case of size 4
-- reg_a = a0_X; reg_b = b3_X; reg_acc = reg_o; Enable sign b; operation : a*b + acc;
"000000100001011000000000100000000001000100001100000011",
--  (1018) multiplication_with_reduction_special_prime_3_16
-- reg_a = a3_X; reg_b = b0_X; reg_acc = reg_o; o3_X = reg_o; Enable sign a; operation : a*b + acc;
"000000100001011000010000100000000000100001100001100011",
--  (1019) multiplication_with_reduction_special_prime_3_17
-- reg_a = a1_X; reg_b = b3_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001011000000000100000100001000100001100100011",
--  (1020) multiplication_with_reduction_special_prime_3_18
-- reg_a = o1_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001011000000000100000000000000100001100110111",
--  (1021) multiplication_with_reduction_special_prime_3_19
-- reg_a = a2_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001011000000000100000000000000100001001000011",
--  (1022) multiplication_with_reduction_special_prime_3_20
-- reg_a = a3_X; reg_b = b1_X; reg_acc = reg_o; Enable sign a; o0_X = reg_o; operation : a*b + acc;
"000000100001011000010000100000000000100100000101100011",
--  (1023) multiplication_with_reduction_special_prime_3_21
-- reg_a = a2_X; reg_b = b3_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001011000000000100000100001000100001101000011",
--  (1024) multiplication_with_reduction_special_prime_3_22
-- reg_a = o2_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001011000000000100000000000000100001101010111",
--  (1025) multiplication_with_reduction_special_prime_3_23
-- reg_a = a3_X; reg_b = b2_X; reg_acc = reg_o; Enable sign a; o1_X = reg_o; operation : a*b + acc;
"000000100001011000010000100000000000101000101001100011",
--  (1026) multiplication_with_reduction_special_prime_3_24
-- reg_a = a3_X; reg_b = b3_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001011000000000100000100001100100001101100011",
--  (1027) multiplication_with_reduction_special_prime_3_25
-- reg_a = o3_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; o3_X = reg_o >> 256; operation : a*b + acc;
"000000100001011001110000100000000000001101001101110111",
--  (1028) multiplication_with_reduction_special_prime_3_26
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (1029) multiplication_with_reduction_special_prime_3_27
-- -- In case of sizes 5, 6, 7, 8
-- reg_a = a0_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001100000011",
--  (1030) multiplication_with_reduction_special_prime_3_28
-- reg_a = a3_X; reg_b = b0_X; reg_acc = reg_o; o3_X = reg_o; operation : a*b + acc;
"000000100001100000010000100000000000010001100001100011",
--  (1031) multiplication_with_reduction_special_prime_3_29
-- reg_a = o0_X; reg_b = primeSP4; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001100000000000100000100000000100010000010111",
--  (1032) multiplication_with_reduction_special_prime_3_30
-- reg_a = a1_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001100100011",
--  (1033) multiplication_with_reduction_special_prime_3_31
-- reg_a = o1_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001100110111",
--  (1034) multiplication_with_reduction_special_prime_3_32
-- reg_a = a2_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001001000011",
--  (1035) multiplication_with_reduction_special_prime_3_33
-- reg_a = a3_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
"001010100001100000000000100000000000000100000101100011",
--  (1036) multiplication_with_reduction_special_prime_3_34
-- In case of size 5
-- reg_a = a0_X; reg_b = b4_X; reg_acc = reg_o; Enable sign b; operation : a*b + acc;
"000000100001100000000000100000000001000100010000000011",
--  (1037) multiplication_with_reduction_special_prime_3_35
-- reg_a = a4_X; reg_b = b0_X; reg_acc = reg_o; o4_X = reg_o; Enable sign a; operation : a*b + acc;
"000000100001100000010000100000000000100010000010000011",
--  (1038) multiplication_with_reduction_special_prime_3_36
-- reg_a = a1_X; reg_b = b4_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001100000000000100000100001000100010000100011",
--  (1039) multiplication_with_reduction_special_prime_3_37
-- reg_a = o1_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100010000110111",
--  (1040) multiplication_with_reduction_special_prime_3_38
-- reg_a = a2_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001101000011",
--  (1041) multiplication_with_reduction_special_prime_3_39
-- reg_a = o2_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001101010111",
--  (1042) multiplication_with_reduction_special_prime_3_40
-- reg_a = a3_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001001100011",
--  (1043) multiplication_with_reduction_special_prime_3_41
-- reg_a = a4_X; reg_b = b1_X; reg_acc = reg_o; o0_X = reg_o; Enable sign a; operation : a*b + acc;
"000000100001100000010000100000000000100100000110000011",
--  (1044) multiplication_with_reduction_special_prime_3_42
-- reg_a = a2_X; reg_b = b4_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001100000000000100000100001000100010001000011",
--  (1045) multiplication_with_reduction_special_prime_3_43
-- reg_a = o2_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100010001010111",
--  (1046) multiplication_with_reduction_special_prime_3_44
-- reg_a = a3_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001101100011",
--  (1047) multiplication_with_reduction_special_prime_3_45
-- reg_a = o3_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001101110111",
--  (1048) multiplication_with_reduction_special_prime_3_46
-- reg_a = a4_X; reg_b = b2_X; reg_acc = reg_o; Enable sign a; o1_X = reg_o; operation : a*b + acc;
"000000100001100000010000100000000000101000101010000011",
--  (1049) multiplication_with_reduction_special_prime_3_47
-- reg_a = a3_X; reg_b = b4_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001100000000000100000100001000100010001100011",
--  (1050) multiplication_with_reduction_special_prime_3_48
-- reg_a = o3_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100010001110111",
--  (1051) multiplication_with_reduction_special_prime_3_49
-- reg_a = a4_X; reg_b = b3_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001100000000000100000000000100100001110000011",
--  (1052) multiplication_with_reduction_special_prime_3_50
-- reg_a = o4_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
"000000100001100000010000100000000000001101001110010111",
--  (1053) multiplication_with_reduction_special_prime_3_51
-- reg_a = a4_X; reg_b = b4_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001100000000000100000100001100100010010000011",
--  (1054) multiplication_with_reduction_special_prime_3_52
-- reg_a = o4_X; reg_b = primeSP4; reg_acc = reg_o; o3_X = reg_o; o4_X = reg_o >> 256; operation : a*b + acc;
"000000100001100001110000100000000000010001110010010111",
--  (1055) multiplication_with_reduction_special_prime_3_53
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (1056) multiplication_with_reduction_special_prime_3_54
-- -- In case of sizes 6, 7, 8
-- reg_a = a0_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010000000011",
--  (1057) multiplication_with_reduction_special_prime_3_55
-- reg_a = a4_X; reg_b = b0_X; reg_acc = reg_o; o4_X = reg_o; operation : a*b + acc;
"000000100001101000010000100000000000010110000010000011",
--  (1058) multiplication_with_reduction_special_prime_3_56
-- reg_a = o0_X; reg_b = primeSP5; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001101000000000100000100000000100010100010111",
--  (1059) multiplication_with_reduction_special_prime_3_57
-- reg_a = a1_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010000100011",
--  (1060) multiplication_with_reduction_special_prime_3_58
-- reg_a = o1_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010000110111",
--  (1061) multiplication_with_reduction_special_prime_3_59
-- reg_a = a2_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001101000011",
--  (1062) multiplication_with_reduction_special_prime_3_60
-- reg_a = o2_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001101010111",
--  (1063) multiplication_with_reduction_special_prime_3_61
-- reg_a = a3_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001001100011",
--  (1064) multiplication_with_reduction_special_prime_3_62
-- reg_a = a4_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
"001111100001101000000000100000000000000100000110000011",
--  (1065) multiplication_with_reduction_special_prime_3_63
-- In case of size 6
-- reg_a = a0_X; reg_b = b5_X; reg_acc = reg_o; Enable sign b; operation : a*b + acc;
"000000100001101000000000100000000001000100010100000011",
--  (1066) multiplication_with_reduction_special_prime_3_64
-- reg_a = a5_X; reg_b = b0_X; reg_acc = reg_o; o5_X = reg_o; Enable sign a; operation : a*b + acc;
"000000100001101000010000100000000000100010100010100011",
--  (1067) multiplication_with_reduction_special_prime_3_65
-- reg_a = a1_X; reg_b = b5_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001101000000000100000100001000100010100100011",
--  (1068) multiplication_with_reduction_special_prime_3_66
-- reg_a = o1_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010100110111",
--  (1069) multiplication_with_reduction_special_prime_3_67
-- reg_a = a2_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010001000011",
--  (1070) multiplication_with_reduction_special_prime_3_68
-- reg_a = o2_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010001010111",
--  (1071) multiplication_with_reduction_special_prime_3_69
-- reg_a = a3_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001101100011",
--  (1072) multiplication_with_reduction_special_prime_3_70
-- reg_a = o3_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001101110111",
--  (1073) multiplication_with_reduction_special_prime_3_71
-- reg_a = a4_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001010000011",
--  (1074) multiplication_with_reduction_special_prime_3_72
-- reg_a = a5_X; reg_b = b1_X; reg_acc = reg_o; o0_X = reg_o; Enable sign a; operation : a*b + acc;
"000000100001101000010000100000000000100100000110100011",
--  (1075) multiplication_with_reduction_special_prime_3_73
-- reg_a = a2_X; reg_b = b5_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001101000000000100000100001000100010101000011",
--  (1076) multiplication_with_reduction_special_prime_3_74
-- reg_a = o2_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010101010111",
--  (1077) multiplication_with_reduction_special_prime_3_75
-- reg_a = a3_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010001100011",
--  (1078) multiplication_with_reduction_special_prime_3_76
-- reg_a = o3_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010001110111",
--  (1079) multiplication_with_reduction_special_prime_3_77
-- reg_a = a4_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001110000011",
--  (1080) multiplication_with_reduction_special_prime_3_78
-- reg_a = o4_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001110010111",
--  (1081) multiplication_with_reduction_special_prime_3_79
-- reg_a = a5_X; reg_b = b2_X; reg_acc = reg_o; Enable sign a; o1_X = reg_o; operation : a*b + acc;
"000000100001101000010000100000000000101000101010100011",
--  (1082) multiplication_with_reduction_special_prime_3_80
-- reg_a = a3_X; reg_b = b5_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001101000000000100000100001000100010101100011",
--  (1083) multiplication_with_reduction_special_prime_3_81
-- reg_a = o3_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010101110111",
--  (1084) multiplication_with_reduction_special_prime_3_82
-- reg_a = a4_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010010000011",
--  (1085) multiplication_with_reduction_special_prime_3_83
-- reg_a = o4_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010010010111",
--  (1086) multiplication_with_reduction_special_prime_3_84
-- reg_a = a5_X; reg_b = b3_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001101000000000100000000000100100001110100011",
--  (1087) multiplication_with_reduction_special_prime_3_85
-- reg_a = o5_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
"000000100001101000010000100000000000001101001110110111",
--  (1088) multiplication_with_reduction_special_prime_3_86
-- reg_a = a4_X; reg_b = b5_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001101000000000100000100001000100010110000011",
--  (1089) multiplication_with_reduction_special_prime_3_87
-- reg_a = o4_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010110010111",
--  (1090) multiplication_with_reduction_special_prime_3_88
-- reg_a = a5_X; reg_b = b4_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001101000000000100000000000100100010010100011",
--  (1091) multiplication_with_reduction_special_prime_3_89
-- reg_a = o5_X; reg_b = primeSP4; reg_acc = reg_o; o3_X = reg_o; operation : a*b + acc;
"000000100001101000010000100000000000010001110010110111",
--  (1092) multiplication_with_reduction_special_prime_3_90
-- reg_a = a5_X; reg_b = b5_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001101000000000100000100001100100010110100011",
--  (1093) multiplication_with_reduction_special_prime_3_91
-- reg_a = o5_X; reg_b = primeSP5; reg_acc = reg_o; o4_X = reg_o; o5_X = reg_o >> 256; operation : a*b + acc;
"000000100001101001110000100000000000010110010110110111",
--  (1094) multiplication_with_reduction_special_prime_3_92
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (1095) multiplication_with_reduction_special_prime_3_93
-- -- In case of sizes 7, 8
-- reg_a = a0_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010100000011",
--  (1096) multiplication_with_reduction_special_prime_3_94
-- reg_a = a5_X; reg_b = b0_X; reg_acc = reg_o; o5_X = reg_o; operation : a*b + acc;
"000000100001110000010000100000000000011010100010100011",
--  (1097) multiplication_with_reduction_special_prime_3_95
-- reg_a = o0_X; reg_b = primeSP6; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001110000000000100000100000000100011000010111",
--  (1098) multiplication_with_reduction_special_prime_3_96
-- reg_a = a1_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010100100011",
--  (1099) multiplication_with_reduction_special_prime_3_97
-- reg_a = o1_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010100110111",
--  (1100) multiplication_with_reduction_special_prime_3_98
-- reg_a = a2_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010001000011",
--  (1101) multiplication_with_reduction_special_prime_3_99
-- reg_a = o2_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010001010111",
--  (1102) multiplication_with_reduction_special_prime_3_100
-- reg_a = a3_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001101100011",
--  (1103) multiplication_with_reduction_special_prime_3_101
-- reg_a = o3_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001101110111",
--  (1104) multiplication_with_reduction_special_prime_3_102
-- reg_a = a4_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001010000011",
--  (1105) multiplication_with_reduction_special_prime_3_103
-- reg_a = a5_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
"010101100001110000000000100000000000000100000110100011",
--  (1106) multiplication_with_reduction_special_prime_3_104
-- -- In case of size 7
-- reg_a = a0_X; reg_b = b6_X; reg_acc = reg_o; Enable sign b; operation : a*b + acc;
"000000100001110000000000100000000001000100011000000011",
--  (1107) multiplication_with_reduction_special_prime_3_105
-- reg_a = a6_X; reg_b = b0_X; reg_acc = reg_o; o6_X = reg_o; Enable sign a; operation : a*b + acc;
"000000100001110000010000100000000000111111000011000011",
--  (1108) multiplication_with_reduction_special_prime_3_106
-- reg_a = a1_X; reg_b = b6_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001110000000000100000100001000100011000100011",
--  (1109) multiplication_with_reduction_special_prime_3_107
-- reg_a = o1_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100011000110111",
--  (1110) multiplication_with_reduction_special_prime_3_108
-- reg_a = a2_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010101000011",
--  (1111) multiplication_with_reduction_special_prime_3_109
-- reg_a = o2_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010101010111",
--  (1112) multiplication_with_reduction_special_prime_3_110
-- reg_a = a3_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010001100011",
--  (1113) multiplication_with_reduction_special_prime_3_111
-- reg_a = o3_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010001110111",
--  (1114) multiplication_with_reduction_special_prime_3_112
-- reg_a = a4_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001110000011",
--  (1115) multiplication_with_reduction_special_prime_3_113
-- reg_a = o4_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001110010111",
--  (1116) multiplication_with_reduction_special_prime_3_114
-- reg_a = a5_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001010100011",
--  (1117) multiplication_with_reduction_special_prime_3_115
-- reg_a = a6_X; reg_b = b1_X; reg_acc = reg_o; o0_X = reg_o; Enable sign a; operation : a*b + acc;
"000000100001110000010000100000000000100100000111000011",
--  (1118) multiplication_with_reduction_special_prime_3_116
-- reg_a = a2_X; reg_b = b6_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001110000000000100000100001000100011001000011",
--  (1119) multiplication_with_reduction_special_prime_3_117
-- reg_a = o2_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100011001010111",
--  (1120) multiplication_with_reduction_special_prime_3_118
-- reg_a = a3_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010101100011",
--  (1121) multiplication_with_reduction_special_prime_3_119
-- reg_a = o3_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010101110111",
--  (1122) multiplication_with_reduction_special_prime_3_120
-- reg_a = a4_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010010000011",
--  (1123) multiplication_with_reduction_special_prime_3_121
-- reg_a = o4_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010010010111",
--  (1124) multiplication_with_reduction_special_prime_3_122
-- reg_a = a5_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001110100011",
--  (1125) multiplication_with_reduction_special_prime_3_123
-- reg_a = o5_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001110110111",
--  (1126) multiplication_with_reduction_special_prime_3_124
-- reg_a = a6_X; reg_b = b2_X; reg_acc = reg_o; o1_X = reg_o; Enable sign a; operation : a*b + acc;
"000000100001110000010000100000000000101000101011000011",
--  (1127) multiplication_with_reduction_special_prime_3_125
-- reg_a = a3_X; reg_b = b6_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001110000000000100000100001000100011001100011",
--  (1128) multiplication_with_reduction_special_prime_3_126
-- reg_a = o3_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100011001110111",
--  (1129) multiplication_with_reduction_special_prime_3_127
-- reg_a = a4_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010110000011",
--  (1130) multiplication_with_reduction_special_prime_3_128
-- reg_a = o4_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010110010111",
--  (1131) multiplication_with_reduction_special_prime_3_129
-- reg_a = a5_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010010100011",
--  (1132) multiplication_with_reduction_special_prime_3_130
-- reg_a = o5_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010010110111",
--  (1133) multiplication_with_reduction_special_prime_3_131
-- reg_a = a6_X; reg_b = b3_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001110000000000100000000000100100001111000011",
--  (1134) multiplication_with_reduction_special_prime_3_132
-- reg_a = o6_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
"000000100001110000010000100000000000001101001111010111",
--  (1135) multiplication_with_reduction_special_prime_3_133
-- reg_a = a4_X; reg_b = b6_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001110000000000100000100001000100011010000011",
--  (1136) multiplication_with_reduction_special_prime_3_134
-- reg_a = o4_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100011010010111",
--  (1137) multiplication_with_reduction_special_prime_3_135
-- reg_a = a5_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010110100011",
--  (1138) multiplication_with_reduction_special_prime_3_136
-- reg_a = o5_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010110110111",
--  (1139) multiplication_with_reduction_special_prime_3_137
-- reg_a = a6_X; reg_b = b4_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001110000000000100000000000100100010011000011",
--  (1140) multiplication_with_reduction_special_prime_3_138
-- reg_a = o6_X; reg_b = primeSP4; reg_acc = reg_o; o3_X = reg_o; operation : a*b + acc;
"000000100001110000010000100000000000010001110011010111",
--  (1141) multiplication_with_reduction_special_prime_3_139
-- reg_a = a5_X; reg_b = b6_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001110000000000100000100001000100011010100011",
--  (1142) multiplication_with_reduction_special_prime_3_140
-- reg_a = o5_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100011010110111",
--  (1143) multiplication_with_reduction_special_prime_3_141
-- reg_a = a6_X; reg_b = b5_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001110000000000100000000000100100010111000011",
--  (1144) multiplication_with_reduction_special_prime_3_142
-- reg_a = o6_X; reg_b = primeSP5; reg_acc = reg_o; o4_X = reg_o; operation : a*b + acc;
"000000100001110000010000100000000000010110010111010111",
--  (1145) multiplication_with_reduction_special_prime_3_143
-- reg_a = a6_X; reg_b = b6_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001110000000000100000100001100100011011000011",
--  (1146) multiplication_with_reduction_special_prime_3_144
-- reg_a = o6_X; reg_b = primeSP6; reg_acc = reg_o; o5_X = reg_o; o6_X = reg_o >> 256; operation : a*b + acc;
"000000100001110001110000100000000000011010111011010111",
--  (1147) multiplication_with_reduction_special_prime_3_145
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (1148) multiplication_with_reduction_special_prime_3_146
-- -- In case of size 8
-- reg_a = a0_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011000000011",
--  (1149) multiplication_with_reduction_special_prime_3_147
-- reg_a = a6_X; reg_b = b0_X; reg_acc = reg_o; o6_X = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000011111000011000011",
--  (1150) multiplication_with_reduction_special_prime_3_148
-- reg_a = o0_X; reg_b = primeSP7; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001111000000000100000100000000100011100010111",
--  (1151) multiplication_with_reduction_special_prime_3_149
-- reg_a = a1_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011000100011",
--  (1152) multiplication_with_reduction_special_prime_3_150
-- reg_a = o1_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011000110111",
--  (1153) multiplication_with_reduction_special_prime_3_151
-- reg_a = a2_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010101000011",
--  (1154) multiplication_with_reduction_special_prime_3_152
-- reg_a = o2_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010101010111",
--  (1155) multiplication_with_reduction_special_prime_3_153
-- reg_a = a3_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010001100011",
--  (1156) multiplication_with_reduction_special_prime_3_154
-- reg_a = o3_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010001110111",
--  (1157) multiplication_with_reduction_special_prime_3_155
-- reg_a = a4_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001110000011",
--  (1158) multiplication_with_reduction_special_prime_3_156
-- reg_a = o4_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001110010111",
--  (1159) multiplication_with_reduction_special_prime_3_157
-- reg_a = a5_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001010100011",
--  (1160) multiplication_with_reduction_special_prime_3_158
-- reg_a = a6_X; reg_b = b1_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100000111000011",
--  (1161) multiplication_with_reduction_special_prime_3_159
-- reg_a = a0_X; reg_b = b7_X; reg_acc = reg_o; Enable sign b; operation : a*b + acc;
"000000100001111000000000100000000001000100011100000011",
--  (1162) multiplication_with_reduction_special_prime_3_160
-- reg_a = a7_X; reg_b = b0_X; reg_acc = reg_o; o7_X = reg_o; Enable sign a; operation : a*b + acc;
"000000100001111000010000100000000000100011100011100011",
--  (1163) multiplication_with_reduction_special_prime_3_161
-- reg_a = a1_X; reg_b = b7_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001111000000000100000100001000100011100100011",
--  (1164) multiplication_with_reduction_special_prime_3_162
-- reg_a = o1_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011100110111",
--  (1165) multiplication_with_reduction_special_prime_3_163
-- reg_a = a2_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011001000011",
--  (1166) multiplication_with_reduction_special_prime_3_164
-- reg_a = o2_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011001010111",
--  (1167) multiplication_with_reduction_special_prime_3_165
-- reg_a = a3_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010101100011",
--  (1168) multiplication_with_reduction_special_prime_3_166
-- reg_a = o3_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010101110111",
--  (1169) multiplication_with_reduction_special_prime_3_167
-- reg_a = a4_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010010000011",
--  (1170) multiplication_with_reduction_special_prime_3_168
-- reg_a = o4_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010010010111",
--  (1171) multiplication_with_reduction_special_prime_3_169
-- reg_a = a5_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001110100011",
--  (1172) multiplication_with_reduction_special_prime_3_170
-- reg_a = o5_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001110110111",
--  (1173) multiplication_with_reduction_special_prime_3_171
-- reg_a = a6_X; reg_b = b2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001011000011",
--  (1174) multiplication_with_reduction_special_prime_3_172
-- reg_a = a7_X; reg_b = b1_X; reg_acc = reg_o; o0_X = reg_o; Enable sign a; operation : a*b + acc;
"000000100001111000010000100000000000100100000111100011",
--  (1175) multiplication_with_reduction_special_prime_3_173
-- reg_a = a2_X; reg_b = b7_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001111000000000100000100001000100011101000011",
--  (1176) multiplication_with_reduction_special_prime_3_174
-- reg_a = o2_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011101010111",
--  (1177) multiplication_with_reduction_special_prime_3_175
-- reg_a = a3_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011001100011",
--  (1178) multiplication_with_reduction_special_prime_3_176
-- reg_a = o3_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011001110111",
--  (1179) multiplication_with_reduction_special_prime_3_177
-- reg_a = a4_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010110000011",
--  (1180) multiplication_with_reduction_special_prime_3_178
-- reg_a = o4_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010110010111",
--  (1181) multiplication_with_reduction_special_prime_3_179
-- reg_a = a5_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010010100011",
--  (1182) multiplication_with_reduction_special_prime_3_180
-- reg_a = o5_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010010110111",
--  (1183) multiplication_with_reduction_special_prime_3_181
-- reg_a = a6_X; reg_b = b3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001111000011",
--  (1184) multiplication_with_reduction_special_prime_3_182
-- reg_a = o6_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001111010111",
--  (1185) multiplication_with_reduction_special_prime_3_183
-- reg_a = a7_X; reg_b = b2_X; reg_acc = reg_o; o1_X = reg_o; Enable sign a; operation : a*b + acc;
"000000100001111000010000100000000000101000101011100011",
--  (1186) multiplication_with_reduction_special_prime_3_184
-- reg_a = a3_X; reg_b = b7_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001111000000000100000100001000100011101100011",
--  (1187) multiplication_with_reduction_special_prime_3_185
-- reg_a = o3_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011101110111",
--  (1188) multiplication_with_reduction_special_prime_3_186
-- reg_a = a4_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011010000011",
--  (1189) multiplication_with_reduction_special_prime_3_187
-- reg_a = o4_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011010010111",
--  (1190) multiplication_with_reduction_special_prime_3_188
-- reg_a = a5_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010110100011",
--  (1191) multiplication_with_reduction_special_prime_3_189
-- reg_a = o5_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010110110111",
--  (1192) multiplication_with_reduction_special_prime_3_190
-- reg_a = a6_X; reg_b = b4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010011000011",
--  (1193) multiplication_with_reduction_special_prime_3_191
-- reg_a = o6_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010011010111",
--  (1194) multiplication_with_reduction_special_prime_3_192
-- reg_a = a7_X; reg_b = b3_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001111000000000100000000000100100001111100011",
--  (1195) multiplication_with_reduction_special_prime_3_193
-- reg_a = o7_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000001101001111110111",
--  (1196) multiplication_with_reduction_special_prime_3_194
-- reg_a = a4_X; reg_b = b7_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001111000000000100000100001000100011110000011",
--  (1197) multiplication_with_reduction_special_prime_3_195
-- reg_a = o4_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011110010111",
--  (1198) multiplication_with_reduction_special_prime_3_196
-- reg_a = a5_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011010100011",
--  (1199) multiplication_with_reduction_special_prime_3_197
-- reg_a = o5_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011010110111",
--  (1200) multiplication_with_reduction_special_prime_3_198
-- reg_a = a6_X; reg_b = b5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010111000011",
--  (1201) multiplication_with_reduction_special_prime_3_199
-- reg_a = o6_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010111010111",
--  (1202) multiplication_with_reduction_special_prime_3_200
-- reg_a = a7_X; reg_b = b4_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001111000000000100000000000100100010011100011",
--  (1203) multiplication_with_reduction_special_prime_3_201
-- reg_a = o7_X; reg_b = primeSP4; reg_acc = reg_o; o3_X = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000010001110011110111",
--  (1204) multiplication_with_reduction_special_prime_3_202
-- reg_a = a5_X; reg_b = b7_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001111000000000100000100001000100011110100011",
--  (1205) multiplication_with_reduction_special_prime_3_203
-- reg_a = o5_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011110110111",
--  (1206) multiplication_with_reduction_special_prime_3_204
-- reg_a = a6_X; reg_b = b6_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011011000011",
--  (1207) multiplication_with_reduction_special_prime_3_205
-- reg_a = o6_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011011010111",
--  (1208) multiplication_with_reduction_special_prime_3_206
-- reg_a = a7_X; reg_b = b5_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001111000000000100000000000100100010111100011",
--  (1209) multiplication_with_reduction_special_prime_3_207
-- reg_a = o7_X; reg_b = primeSP5; reg_acc = reg_o; o4_X = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000010110010111110111",
--  (1210) multiplication_with_reduction_special_prime_3_208
-- reg_a = a6_X; reg_b = b7_X; reg_acc = reg_o >> 256; Enable sign b; operation : a*b + acc;
"000000100001111000000000100000100001000100011111000011",
--  (1211) multiplication_with_reduction_special_prime_3_209
-- reg_a = o6_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011111010111",
--  (1212) multiplication_with_reduction_special_prime_3_210
-- reg_a = a7_X; reg_b = b6_X; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
"000000100001111000000000100000000000100100011011100011",
--  (1213) multiplication_with_reduction_special_prime_3_211
-- reg_a = o7_X; reg_b = primeSP6; reg_acc = reg_o; o5_X = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000011010111011110111",
--  (1214) multiplication_with_reduction_special_prime_3_212
-- reg_a = a7_X; reg_b = b7_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001111000000000100000100001100100011111100011",
--  (1215) multiplication_with_reduction_special_prime_3_213
-- reg_a = o7_X; reg_b = primeSP7; reg_acc = reg_o; o6_X = reg_o; o7_X = reg_o >> 256; operation : a*b + acc;
"000000100001111001110000100000000000011111011111110111",
--  (1216) multiplication_with_reduction_special_prime_3_214
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (1217) square_with_reduction_0
-- -- In case of size 1
-- reg_a = a0_X; reg_b = a0_X; reg_acc = 0; Enable sign a,b; operation : a*b + acc;
"000000100001000000000000100000010001100100000000000011",
--  (1218) square_with_reduction_1
-- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o0_X = reg_y; operation : keep accumulator;
"000000100001000000011000110000000100000100000000011011",
--  (1219) square_with_reduction_2
-- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
"000000100001000000000000100000000010000100000000010011",
--  (1220) square_with_reduction_3
-- reg_a = 0; reg_b = 0; reg_acc = reg_o >> 256; o0_X = reg_o; operation : a*b + acc;
"000000100001000000010000100000101110000100000000000011",
--  (1221) square_with_reduction_4
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (1222) square_with_reduction_5
-- -- In case of 2, 3, 4, 5, 6, 7, 8
-- reg_a = a0_X; reg_b = a0_X; reg_acc = 0; operation : a*b + acc;
"000000100001001000000000100000010000000100000000000011",
--  (1223) square_with_reduction_6
-- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o0_X = reg_y; operation : keep accumulator;
"000000100001001000011000110000000100000100000000011011",
--  (1224) square_with_reduction_7
-- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
"000000100001001000000000100000000010000100000000010011",
--  (1225) square_with_reduction_8
-- reg_a = o0_X; reg_b = prime1; reg_acc = reg_o >> 256; operation : a*b + acc;
"000011100001001000000000100000100000000100000100010111",
--  (1226) square_with_reduction_9
-- -- In case of size 2
-- reg_a = a0_X; reg_b = a1_X; reg_acc = reg_o; Enable sign b; operation : 2*a*b + acc;
"000000100001001000000100100000000001000100000100000011",
--  (1227) square_with_reduction_10
-- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o1_X = reg_y; operation : keep accumulator;
"000000100001001000011000110000000100001000100000111011",
--  (1228) square_with_reduction_11
-- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
"000000100001001000000000100000000010000100000000110011",
--  (1229) square_with_reduction_12
-- reg_a = a1_X; reg_b = a1_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001001000000000100000100001100100000100100011",
--  (1230) square_with_reduction_13
-- reg_a = o1_X; reg_b = prime1; reg_acc = reg_o; o0_X = reg_o; o1_X = reg_o >> 256; operation : a*b + acc;
"000000100001001001110000100000000000000100000100110111",
--  (1231) square_with_reduction_14
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (1232) square_with_reduction_15
-- -- Others cases
-- reg_a = a0_X; reg_b = a1_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001010000000100100000000000000100000100000011",
--  (1233) square_with_reduction_16
-- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o1_X = reg_y; operation : keep accumulator;
"000000100001010000011000110000000100001000100000011011",
--  (1234) square_with_reduction_17
-- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
"000000100001010000000000100000000010000100000000010011",
--  (1235) square_with_reduction_18
-- reg_a = o0_X; reg_b = prime2; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001010000000000100000100000000100001000010111",
--  (1236) square_with_reduction_19
-- reg_a = a1_X; reg_b = a1_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001010000000000100000000000000100000100100011",
--  (1237) square_with_reduction_20
-- reg_a = o1_X; reg_b = prime1; reg_acc = reg_o; operation : a*b + acc;
"000101000001010000000000100000000000000100000100110111",
--  (1238) square_with_reduction_21
-- -- In case of size 3
-- reg_a = a0_X; reg_b = a2_X; reg_acc = reg_o; Enable sign b; operation : 2*a*b + acc;
"000000100001010000000100100000000001000100001000000011",
--  (1239) square_with_reduction_22
-- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o2_X = reg_y; operation : keep accumulator;
"000000100001010000011000110000000100001101000000011011",
--  (1240) square_with_reduction_23
-- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
"000000100001010000000000100000000010000100000000010011",
--  (1241) square_with_reduction_24
-- reg_a = a1_X; reg_b = a2_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001010000000100100000100001000100001000100011",
--  (1242) square_with_reduction_25
-- reg_a = o1_X; reg_b = prime2; reg_acc = reg_o; operation : a*b + acc;
"000000100001010000000000100000000000000100001000110111",
--  (1243) square_with_reduction_26
-- reg_a = o2_X; reg_b = prime1; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
"000000100001010000010000100000000000000100000101010111",
--  (1244) square_with_reduction_27
-- reg_a = a2_X; reg_b = a2_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001010000000000100000100001100100001001000011",
--  (1245) square_with_reduction_28
-- reg_a = o2_X; reg_b = prime2; reg_acc = reg_o; o1_X = reg_o; o2_X = reg_o >> 256; operation : a*b + acc;
"000000100001010001110000100000000000001000101001010111",
--  (1246) square_with_reduction_29
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (1247) square_with_reduction_30
-- -- Other cases
-- reg_a = a0_X; reg_b = a2_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001011000000100100000000000000100001000000011",
--  (1248) square_with_reduction_31
-- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o2_X = reg_y; operation : keep accumulator;
"000000100001011000011000110000000100001101000000011011",
--  (1249) square_with_reduction_32
-- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
"000000100001011000000000100000000010000100000000010011",
--  (1250) square_with_reduction_33
-- reg_a = o0_X; reg_b = prime3; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001011000000000100000100000000100001100010111",
--  (1251) square_with_reduction_34
-- reg_a = a1_X; reg_b = a2_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001011000000100100000000000000100001000100011",
--  (1252) square_with_reduction_35
-- reg_a = o1_X; reg_b = prime2; reg_acc = reg_o; operation : a*b + acc;
"000000100001011000000000100000000000000100001000110111",
--  (1253) square_with_reduction_36
-- reg_a = o2_X; reg_b = prime1; reg_acc = reg_o; operation : a*b + acc;
"000111100001011000000000100000000000000100000101010111",
--  (1254) square_with_reduction_37
-- In case of size 4
-- reg_a = a0_X; reg_b = a3_X; reg_acc = reg_o; Enable sign b; operation : 2*a*b + acc;
"000000100001011000000100100000000001000100001100000011",
--  (1255) square_with_reduction_38
-- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o3_X = reg_y; operation : keep accumulator;
"000000100001011000011000110000000100010001100000011011",
--  (1256) square_with_reduction_39
-- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
"000000100001011000000000100000000010000100000000010011",
--  (1257) square_with_reduction_40
-- reg_a = a1_X; reg_b = a3_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001011000000100100000100001000100001100100011",
--  (1258) square_with_reduction_41
-- reg_a = o1_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
"000000100001011000000000100000000000000100001100110111",
--  (1259) square_with_reduction_42
-- reg_a = a2_X; reg_b = a2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001011000000000100000000000000100001001000011",
--  (1260) square_with_reduction_43
-- reg_a = o2_X; reg_b = prime2; reg_acc = reg_o; operation : a*b + acc;
"000000100001011000000000100000000000000100001001010111",
--  (1261) square_with_reduction_44
-- reg_a = o3_X; reg_b = prime1; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
"000000100001011000010000100000000000000100000101110111",
--  (1262) square_with_reduction_45
-- reg_a = a2_X; reg_b = a3_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001011000000100100000100001000100001101000011",
--  (1263) square_with_reduction_46
-- reg_a = o2_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
"000000100001011000000000100000000000000100001101010111",
--  (1264) square_with_reduction_47
-- reg_a = o3_X; reg_b = prime2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
"000000100001011000010000100000000000001000101001110111",
--  (1265) square_with_reduction_48
-- reg_a = a3_X; reg_b = a3_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001011000000000100000100001100100001101100011",
--  (1266) square_with_reduction_49
-- reg_a = o3_X; reg_b = prime3; reg_acc = reg_o; o2_X = reg_o; o3_X = reg_o >> 256; operation : a*b + acc;
"000000100001011001110000100000000000001101001101110111",
--  (1267) square_with_reduction_50
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (1268) square_with_reduction_51
-- -- Other cases
-- reg_a = a0_X; reg_b = a3_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001100000000100100000000000000100001100000011",
--  (1269) square_with_reduction_52
-- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o3_X = reg_y; operation : keep accumulator;
"000000100001100000011000110000000100010001100000011011",
--  (1270) square_with_reduction_53
-- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000010000100000000010011",
--  (1271) square_with_reduction_54
-- reg_a = o0_X; reg_b = prime4; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001100000000000100000100000000100010000010111",
--  (1272) square_with_reduction_55
-- reg_a = a1_X; reg_b = a3_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001100000000100100000000000000100001100100011",
--  (1273) square_with_reduction_56
-- reg_a = o1_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001100110111",
--  (1274) square_with_reduction_57
-- reg_a = a2_X; reg_b = a2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001001000011",
--  (1275) square_with_reduction_58
-- reg_a = o2_X; reg_b = prime2; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001001010111",
--  (1276) square_with_reduction_59
-- reg_a = o3_X; reg_b = prime1; reg_acc = reg_o; operation : a*b + acc;
"001010100001100000000000100000000000000100000101110111",
--  (1277) square_with_reduction_60
-- -- In case of size 5
-- reg_a = a0_X; reg_b = a4_X; reg_acc = reg_o; Enable sign b; operation : 2*a*b + acc;
"000000100001100000000100100000000001000100010000000011",
--  (1278) square_with_reduction_61
-- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o4_X = reg_y; operation : keep accumulator;
"000000100001100000011000110000000100010110000000011011",
--  (1279) square_with_reduction_62
-- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000010000100000000010011",
--  (1280) square_with_reduction_63
-- reg_a = a1_X; reg_b = a4_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001100000000100100000100001000100010000100011",
--  (1281) square_with_reduction_64
-- reg_a = o1_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100010000110111",
--  (1282) square_with_reduction_65
-- reg_a = a2_X; reg_b = a3_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001100000000100100000000000000100001101000011",
--  (1283) square_with_reduction_66
-- reg_a = o2_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001101010111",
--  (1284) square_with_reduction_67
-- reg_a = o3_X; reg_b = prime2; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001001110111",
--  (1285) square_with_reduction_68
-- reg_a = o4_X; reg_b = prime1; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
"000000100001100000010000100000000000000100000110010111",
--  (1286) square_with_reduction_69
-- reg_a = a2_X; reg_b = a4_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001100000000100100000100001000100010001000011",
--  (1287) square_with_reduction_70
-- reg_a = o2_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100010001010111",
--  (1288) square_with_reduction_71
-- reg_a = a3_X; reg_b = a3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001101100011",
--  (1289) square_with_reduction_72
-- reg_a = o3_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001101110111",
--  (1290) square_with_reduction_73
-- reg_a = o4_X; reg_b = prime2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
"000000100001100000010000100000000000001000101010010111",
--  (1291) square_with_reduction_74
-- reg_a = a3_X; reg_b = a4_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001100000000100100000100001000100010001100011",
--  (1292) square_with_reduction_75
-- reg_a = o3_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100010001110111",
--  (1293) square_with_reduction_76
-- reg_a = o4_X; reg_b = prime3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
"000000100001100000010000100000000000001101001110010111",
--  (1294) square_with_reduction_77
-- reg_a = a4_X; reg_b = a4_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001100000000000100000100001100100010010000011",
--  (1295) square_with_reduction_78
-- reg_a = o4_X; reg_b = prime4; reg_acc = reg_o; o3_X = reg_o; o4_X = reg_o >> 256; operation : a*b + acc;
"000000100001100001110000100000000000010001110010010111",
--  (1296) square_with_reduction_79
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (1297) square_with_reduction_80
-- -- Other cases
-- reg_a = a0_X; reg_b = a4_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001101000000100100000000000000100010000000011",
--  (1298) square_with_reduction_81
-- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o4_X = reg_y; operation : keep accumulator;
"000000100001101000011000110000000100010110000000011011",
--  (1299) square_with_reduction_82
-- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000010000100000000010011",
--  (1300) square_with_reduction_83
-- reg_a = o0_X; reg_b = prime5; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001101000000000100000100000000100010100010111",
--  (1301) square_with_reduction_84
-- reg_a = a1_X; reg_b = a4_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001101000000100100000000000000100010000100011",
--  (1302) square_with_reduction_85
-- reg_a = o1_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010000110111",
--  (1303) square_with_reduction_86
-- reg_a = a2_X; reg_b = a3_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001101000000100100000000000000100001101000011",
--  (1304) square_with_reduction_87
-- reg_a = o2_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001101010111",
--  (1305) square_with_reduction_88
-- reg_a = o3_X; reg_b = prime2; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001001110111",
--  (1306) square_with_reduction_89
-- reg_a = o4_X; reg_b = prime1; reg_acc = reg_o; operation : a*b + acc;
"001110100001101000000000100000000000000100000110010111",
--  (1307) square_with_reduction_90
-- -- In case of size 6
-- reg_a = a0_X; reg_b = a5_X; reg_acc = reg_o; Enable sign b; operation : 2*a*b + acc;
"000000100001101000000100100000000001000100010100000011",
--  (1308) square_with_reduction_91
-- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o5_X = reg_y; operation : keep accumulator;
"000000100001101000011000110000000100011010100000011011",
--  (1309) square_with_reduction_92
-- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000010000100000000010011",
--  (1310) square_with_reduction_93
-- reg_a = a1_X; reg_b = a5_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001101000000100100000100001000100010100100011",
--  (1311) square_with_reduction_94
-- reg_a = o1_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010100110111",
--  (1312) square_with_reduction_95
-- reg_a = a2_X; reg_b = a4_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001101000000100100000000000000100010001000011",
--  (1313) square_with_reduction_96
-- reg_a = o2_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010001010111",
--  (1314) square_with_reduction_97
-- reg_a = a3_X; reg_b = a3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001101100011",
--  (1315) square_with_reduction_98
-- reg_a = o3_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001101110111",
--  (1316) square_with_reduction_99
-- reg_a = o4_X; reg_b = prime2; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001010010111",
--  (1317) square_with_reduction_100
-- reg_a = o5_X; reg_b = prime1; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
"000000100001101000010000100000000000000100000110110111",
--  (1318) square_with_reduction_101
-- reg_a = a2_X; reg_b = a5_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001101000000100100000100001000100010101000011",
--  (1319) square_with_reduction_102
-- reg_a = o2_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010101010111",
--  (1320) square_with_reduction_103
-- reg_a = a3_X; reg_b = a4_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001101000000100100000000000000100010001100011",
--  (1321) square_with_reduction_104
-- reg_a = o3_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010001110111",
--  (1322) square_with_reduction_105
-- reg_a = o4_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001110010111",
--  (1323) square_with_reduction_106
-- reg_a = o5_X; reg_b = prime2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
"000000100001101000010000100000000000001000101010110111",
--  (1324) square_with_reduction_107
-- reg_a = a3_X; reg_b = a5_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001101000000100100000100001000100010101100011",
--  (1325) square_with_reduction_108
-- reg_a = o3_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010101110111",
--  (1326) square_with_reduction_109
-- reg_a = a4_X; reg_b = a4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010010000011",
--  (1327) square_with_reduction_110
-- reg_a = o4_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010010010111",
--  (1328) square_with_reduction_111
-- reg_a = o5_X; reg_b = prime3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
"000000100001101000010000100000000000001101001110110111",
--  (1329) square_with_reduction_112
-- reg_a = a4_X; reg_b = a5_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001101000000100100000100001000100010110000011",
--  (1330) square_with_reduction_113
-- reg_a = o4_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010110010111",
--  (1331) square_with_reduction_114
-- reg_a = o5_X; reg_b = prime4; reg_acc = reg_o; o3_X = reg_o; operation : a*b + acc;
"000000100001101000010000100000000000010001110010110111",
--  (1332) square_with_reduction_115
-- reg_a = a5_X; reg_b = a5_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001101000000000100000100001100100010110100011",
--  (1333) square_with_reduction_116
-- reg_a = o5_X; reg_b = prime5; reg_acc = reg_o; o4_X = reg_o; o5_X = reg_o >> 256; operation : a*b + acc;
"000000100001101001110000100000000000010110010110110111",
--  (1334) square_with_reduction_117
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (1335) square_with_reduction_118
-- -- Other cases
-- reg_a = a0_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001110000000100100000000000000100010100000011",
--  (1336) square_with_reduction_119
-- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o5_X = reg_y; operation : keep accumulator;
"000000100001110000011000110000000100010110100000011011",
--  (1337) square_with_reduction_120
-- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000010000100000000010011",
--  (1338) square_with_reduction_121
-- reg_a = o0_X; reg_b = prime6; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001110000000000100000100000000100011000010111",
--  (1339) square_with_reduction_122
-- reg_a = a1_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001110000000100100000000000000100010100100011",
--  (1340) square_with_reduction_123
-- reg_a = o1_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010100110111",
--  (1341) square_with_reduction_124
-- reg_a = a2_X; reg_b = a4_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001110000000100100000000000000100010001000011",
--  (1342) square_with_reduction_125
-- reg_a = o2_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010001010111",
--  (1343) square_with_reduction_126
-- reg_a = a3_X; reg_b = a3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001101100011",
--  (1344) square_with_reduction_127
-- reg_a = o3_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001101110111",
--  (1345) square_with_reduction_128
-- reg_a = o4_X; reg_b = prime2; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001010010111",
--  (1346) square_with_reduction_129
-- reg_a = o5_X; reg_b = prime1; reg_acc = reg_o; operation : a*b + acc;
"010011000001110000000000100000000000000100000110110111",
--  (1347) square_with_reduction_130
-- -- In case of size 7
-- reg_a = a0_X; reg_b = a6_X; reg_acc = reg_o; Enable sign b; operation : 2*a*b + acc;
"000000100001110000000100100000000001000100011000000011",
--  (1348) square_with_reduction_131
-- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o6_X = reg_y; operation : keep accumulator;
"000000100001110000011000110000000100011111000000011011",
--  (1349) square_with_reduction_132
-- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000010000100000000010011",
--  (1350) square_with_reduction_133
-- reg_a = a1_X; reg_b = a6_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001110000000100100000100001000100011000100011",
--  (1351) square_with_reduction_134
-- reg_a = o1_X; reg_b = prime6; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100011000110111",
--  (1352) square_with_reduction_135
-- reg_a = a2_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001110000000100100000000000000100010101000011",
--  (1353) square_with_reduction_136
-- reg_a = o2_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010101010111",
--  (1354) square_with_reduction_137
-- reg_a = a3_X; reg_b = a4_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001110000000100100000000000000100010001100011",
--  (1355) square_with_reduction_138
-- reg_a = o3_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010001110111",
--  (1356) square_with_reduction_139
-- reg_a = o4_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001110010111",
--  (1357) square_with_reduction_140
-- reg_a = o5_X; reg_b = prime2; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001010110111",
--  (1358) square_with_reduction_141
-- reg_a = o6_X; reg_b = prime1; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
"000000100001110000010000100000000000000100000111010111",
--  (1359) square_with_reduction_142
-- reg_a = a2_X; reg_b = a6_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001110000000100100000100001000100011001000011",
--  (1360) square_with_reduction_143
-- reg_a = o2_X; reg_b = prime6; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100011001010111",
--  (1361) square_with_reduction_144
-- reg_a = a3_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001110000000100100000000000000100010101100011",
--  (1362) square_with_reduction_145
-- reg_a = o3_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010101110111",
--  (1363) square_with_reduction_146
-- reg_a = a4_X; reg_b = a4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010010000011",
--  (1364) square_with_reduction_147
-- reg_a = o4_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010010010111",
--  (1365) square_with_reduction_148
-- reg_a = o5_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001110110111",
--  (1366) square_with_reduction_149
-- reg_a = o6_X; reg_b = prime2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
"000000100001110000010000100000000000001000101011010111",
--  (1367) square_with_reduction_150
-- reg_a = a3_X; reg_b = a6_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001110000000100100000100001000100011001100011",
--  (1368) square_with_reduction_151
-- reg_a = o3_X; reg_b = prime6; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100011001110111",
--  (1369) square_with_reduction_152
-- reg_a = a4_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001110000000100100000000000000100010110000011",
--  (1370) square_with_reduction_153
-- reg_a = o4_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010110010111",
--  (1371) square_with_reduction_154
-- reg_a = o5_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010010110111",
--  (1372) square_with_reduction_155
-- reg_a = o6_X; reg_b = prime3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
"000000100001110000010000100000000000001101001111010111",
--  (1373) square_with_reduction_156
-- reg_a = a4_X; reg_b = a6_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001110000000100100000100001000100011010000011",
--  (1374) square_with_reduction_157
-- reg_a = o4_X; reg_b = prime6; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100011010010111",
--  (1375) square_with_reduction_158
-- reg_a = a5_X; reg_b = a5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010110100011",
--  (1376) square_with_reduction_159
-- reg_a = o5_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010110110111",
--  (1377) square_with_reduction_160
-- reg_a = o6_X; reg_b = prime4; reg_acc = reg_o; o3_X = reg_o; operation : a*b + acc;
"000000100001110000010000100000000000010001110011010111",
--  (1378) square_with_reduction_161
-- reg_a = a5_X; reg_b = a6_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001110000000100100000100001000100011010100011",
--  (1379) square_with_reduction_162
-- reg_a = o5_X; reg_b = prime6; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100011010110111",
--  (1380) square_with_reduction_163
-- reg_a = o6_X; reg_b = prime5; reg_acc = reg_o; o4_X = reg_o; operation : a*b + acc;
"000000100001110000010000100000000000010110010111010111",
--  (1381) square_with_reduction_164
-- reg_a = a6_X; reg_b = a6_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001110000000000100000100001100100011011000011",
--  (1382) square_with_reduction_165
-- reg_a = o6_X; reg_b = prime6; reg_acc = reg_o; o5_X = reg_o; o6_X = reg_o >> 256; operation : a*b + acc;
"000000100001110001110000100000000000011010111011010111",
--  (1383) square_with_reduction_166
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (1384) square_with_reduction_167
-- -- In case of size 8
-- reg_a = a0_X; reg_b = a6_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001111000000100100000000000000100011000000011",
--  (1385) square_with_reduction_168
-- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o6_X = reg_y; operation : keep accumulator;
"000000100001111000011000110000000100011111000000011011",
--  (1386) square_with_reduction_169
-- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000010000100000000010011",
--  (1387) square_with_reduction_170
-- reg_a = o0_X; reg_b = prime7; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001111000000000100000100000000100011100010111",
--  (1388) square_with_reduction_171
-- reg_a = a1_X; reg_b = a6_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001111000000100100000000000000100011000100011",
--  (1389) square_with_reduction_172
-- reg_a = o1_X; reg_b = prime6; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011000110111",
--  (1390) square_with_reduction_173
-- reg_a = a2_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001111000000100100000000000000100010101000011",
--  (1391) square_with_reduction_174
-- reg_a = o2_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010101010111",
--  (1392) square_with_reduction_175
-- reg_a = a3_X; reg_b = a4_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001111000000100100000000000000100010001100011",
--  (1393) square_with_reduction_176
-- reg_a = o3_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010001110111",
--  (1394) square_with_reduction_177
-- reg_a = o4_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001010010111",
--  (1395) square_with_reduction_178
-- reg_a = o5_X; reg_b = prime2; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001010110111",
--  (1396) square_with_reduction_179
-- reg_a = o6_X; reg_b = prime1; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100000111010111",
--  (1397) square_with_reduction_180
-- reg_a = a0_X; reg_b = a7_X; reg_acc = reg_o; Enable sign b; operation : 2*a*b + acc;
"000000100001111000000100100000000001000100011100000011",
--  (1398) square_with_reduction_181
-- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o7_X = reg_y; operation : keep accumulator;
"000000100001111000011000110000000100000011100000011011",
--  (1399) square_with_reduction_182
-- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000010000100000000010011",
--  (1400) square_with_reduction_183
-- reg_a = a1_X; reg_b = a7_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001111000000100100000100001000100011100100011",
--  (1401) square_with_reduction_184
-- reg_a = o1_X; reg_b = prime7; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011100110111",
--  (1402) square_with_reduction_185
-- reg_a = a2_X; reg_b = a6_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001111000000100100000000000000100011001000011",
--  (1403) square_with_reduction_186
-- reg_a = o2_X; reg_b = prime6; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011001010111",
--  (1404) square_with_reduction_187
-- reg_a = a3_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001111000000100100000000000000100010101100011",
--  (1405) square_with_reduction_188
-- reg_a = o3_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010101110111",
--  (1406) square_with_reduction_189
-- reg_a = a4_X; reg_b = a4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010010000011",
--  (1407) square_with_reduction_190
-- reg_a = o4_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010010010111",
--  (1408) square_with_reduction_191
-- reg_a = o5_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001110110111",
--  (1409) square_with_reduction_192
-- reg_a = o6_X; reg_b = prime2; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001011010111",
--  (1410) square_with_reduction_193
-- reg_a = o7_X; reg_b = prime1; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000000100000111110111",
--  (1411) square_with_reduction_194
-- reg_a = a2_X; reg_b = a7_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001111000000100100000100001000100011101000011",
--  (1412) square_with_reduction_195
-- reg_a = o2_X; reg_b = prime7; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011101010111",
--  (1413) square_with_reduction_196
-- reg_a = a3_X; reg_b = a6_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001111000000100100000000000000100011001100011",
--  (1414) square_with_reduction_197
-- reg_a = o3_X; reg_b = prime6; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011001110111",
--  (1415) square_with_reduction_198
-- reg_a = a4_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001111000000100100000000000000100010110000011",
--  (1416) square_with_reduction_199
-- reg_a = o4_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010110010111",
--  (1417) square_with_reduction_200
-- reg_a = o5_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010010110111",
--  (1418) square_with_reduction_201
-- reg_a = o6_X; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001111010111",
--  (1419) square_with_reduction_202
-- reg_a = o7_X; reg_b = prime2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000001000101011110111",
--  (1420) square_with_reduction_203
-- reg_a = a3_X; reg_b = a7_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001111000000100100000100001000100011101100011",
--  (1421) square_with_reduction_204
-- reg_a = o3_X; reg_b = prime7; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011101110111",
--  (1422) square_with_reduction_205
-- reg_a = a4_X; reg_b = a6_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001111000000100100000000000000100011010000011",
--  (1423) square_with_reduction_206
-- reg_a = o4_X; reg_b = prime6; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011010010111",
--  (1424) square_with_reduction_207
-- reg_a = a5_X; reg_b = a5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010110100011",
--  (1425) square_with_reduction_208
-- reg_a = o5_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010110110111",
--  (1426) square_with_reduction_209
-- reg_a = o6_X; reg_b = prime4; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010011010111",
--  (1427) square_with_reduction_210
-- reg_a = o7_X; reg_b = prime3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000001101001111110111",
--  (1428) square_with_reduction_211
-- reg_a = a4_X; reg_b = a7_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001111000000100100000100001000100011110000011",
--  (1429) square_with_reduction_212
-- reg_a = o4_X; reg_b = prime7; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011110010111",
--  (1430) square_with_reduction_213
-- reg_a = a5_X; reg_b = a6_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001111000000100100000000000000100011010100011",
--  (1431) square_with_reduction_214
-- reg_a = o5_X; reg_b = prime6; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011010110111",
--  (1432) square_with_reduction_215
-- reg_a = o6_X; reg_b = prime5; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010111010111",
--  (1433) square_with_reduction_216
-- reg_a = o7_X; reg_b = prime4; reg_acc = reg_o; o3_X = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000010001110011110111",
--  (1434) square_with_reduction_217
-- reg_a = a5_X; reg_b = a7_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001111000000100100000100001000100011110100011",
--  (1435) square_with_reduction_218
-- reg_a = o5_X; reg_b = prime7; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011110110111",
--  (1436) square_with_reduction_219
-- reg_a = a6_X; reg_b = a6_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011011000011",
--  (1437) square_with_reduction_220
-- reg_a = o6_X; reg_b = prime6; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011011010111",
--  (1438) square_with_reduction_221
-- reg_a = o7_X; reg_b = prime5; reg_acc = reg_o; o4_X = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000010110010111110111",
--  (1439) square_with_reduction_222
-- reg_a = a6_X; reg_b = a7_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001111000000100100000100001000100011111000011",
--  (1440) square_with_reduction_223
-- reg_a = o6_X; reg_b = prime7; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011111010111",
--  (1441) square_with_reduction_224
-- reg_a = o7_X; reg_b = prime6; reg_acc = reg_o; o5_X = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000011010111011110111",
--  (1442) square_with_reduction_225
-- reg_a = a7_X; reg_b = a7_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001111000000000100000100001100100011111100011",
--  (1443) square_with_reduction_226
-- reg_a = o7_X; reg_b = prime7; reg_acc = reg_o; o6_X = reg_o; o7_X = reg_o >> 256; operation : a*b + acc;
"000000100001111001110000100000000000011111011111110111",
--  (1444) square_with_reduction_227
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (1445) square_with_reduction_special_prime_1_0
-- -- In case of size 1
-- reg_a = a0_X; reg_b = a0_X; reg_acc = 0; Enable sign a,b; operation : a*b + acc;
"000000100001000000000000100000010001100100000000000011",
--  (1446) square_with_reduction_special_prime_1_1
-- reg_a = 0; reg_b = 0; reg_acc = reg_o >> 256; o0_X = reg_o; operation : a*b + acc;
"000000100001000000010000100000101110000100000000000011",
--  (1447) square_with_reduction_special_prime_1_2
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (1448) square_with_reduction_special_prime_1_3
-- -- In case of size 2, 3, 4, 5, 6, 7, 8
-- reg_a = a0_X; reg_b = a0_X; reg_acc = 0; o0_X = reg_o; operation : a*b + acc;
"000000100001001000010000100000010000000100000000000011",
--  (1449) square_with_reduction_special_prime_1_4
-- reg_a = reg_o; reg_b = primeSP1; reg_acc = reg_o >> 256; operation : a*b + acc;
"000010100001001000000000100000100100001000100100010111",
--  (1450) square_with_reduction_special_prime_1_5
-- -- In case of size 2
-- reg_a = a0_X; reg_b = a1_X; reg_acc = reg_o; o1_X = reg_o; Enable sign b; operation : 2*a*b + acc;
"000000100001001000010100100000000001001000100100000011",
--  (1451) square_with_reduction_special_prime_1_6
-- reg_a = a1_X; reg_b = a1_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001001000000000100000100001100100000100100011",
--  (1452) square_with_reduction_special_prime_1_7
-- reg_a = o1_X; reg_b = primeSP1; reg_acc = reg_o; o0_X = reg_o; o1_X = reg_o >> 256; operation : a*b + acc;
"000000100001001001110000100000000000000100000100110111",
--  (1453) square_with_reduction_special_prime_1_8
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (1454) square_with_reduction_special_prime_1_9
-- -- In case of size 3, 4, 5, 6, 7, 8
-- reg_a = a0_X; reg_b = a1_X; reg_acc = reg_o; o1_X = reg_o; operation : 2*a*b + acc;
"000000100001010000010100100000000000001000100100000011",
--  (1455) square_with_reduction_special_prime_1_10
-- reg_a = o0_X; reg_b = primeSP2; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001010000000000100000100000000100001000010111",
--  (1456) square_with_reduction_special_prime_1_11
-- reg_a = a1_X; reg_b = a1_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001010000000000100000000000000100000100100011",
--  (1457) square_with_reduction_special_prime_1_12
-- reg_a = o1_X; reg_b = primeSP1; reg_acc = reg_o; operation : a*b + acc;
"000100000001010000000000100000000000001101000100110111",
--  (1458) square_with_reduction_special_prime_1_13
-- -- In case of size 3
-- reg_a = a0_X; reg_b = a2_X; reg_acc = reg_o; o2_X = reg_o; Enable sign b; operation : 2*a*b + acc;
"000000100001010000010100100000000001001101001000000011",
--  (1459) square_with_reduction_special_prime_1_14
-- reg_a = a1_X; reg_b = a2_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001010000000100100000100001000100001000100011",
--  (1460) square_with_reduction_special_prime_1_15
-- reg_a = o1_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
"000000100001010000000000100000000000000100001000110111",
--  (1461) square_with_reduction_special_prime_1_16
-- reg_a = o2_X; reg_b = primeSP1; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
"000000100001010000010000100000000000000100000101010111",
--  (1462) square_with_reduction_special_prime_1_17
-- reg_a = a2_X; reg_b = a2_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001010000000000100000100001100100001001000011",
--  (1463) square_with_reduction_special_prime_1_18
-- reg_a = o2_X; reg_b = primeSP2; reg_acc = reg_o; o1_X = reg_o; o2_X = reg_o >> 256; operation : a*b + acc;
"000000100001010001110000100000000000001000101001010111",
--  (1464) square_with_reduction_special_prime_1_19
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (1465) square_with_reduction_special_prime_1_20
-- -- In case of sizes 4, 5, 6, 7, 8
-- reg_a = a0_X; reg_b = a2_X; reg_acc = reg_o; o2_X = reg_o; operation : 2*a*b + acc;
"000000100001011000010100100000000000001101001000000011",
--  (1466) square_with_reduction_special_prime_1_21
-- reg_a = o0_X; reg_b = primeSP3; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001011000000000100000100000000100001100010111",
--  (1467) square_with_reduction_special_prime_1_22
-- reg_a = a1_X; reg_b = a2_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001011000000100100000000000000100001000100011",
--  (1468) square_with_reduction_special_prime_1_23
-- reg_a = o1_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
"000000100001011000000000100000000000000100001000110111",
--  (1469) square_with_reduction_special_prime_1_24
-- reg_a = o2_X; reg_b = primeSP1; reg_acc = reg_o; operation : a*b + acc;
"000110100001011000000000100000000000000100000101010111",
--  (1470) square_with_reduction_special_prime_1_25
-- -- In case of size 4
-- reg_a = a0_X; reg_b = a3_X; reg_acc = reg_o; o3_X = reg_o; Enable sign b; operation : 2*a*b + acc;
"000000100001011000010100100000000001010001101100000011",
--  (1471) square_with_reduction_special_prime_1_26
-- reg_a = a1_X; reg_b = a3_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001011000000100100000100001000100001100100011",
--  (1472) square_with_reduction_special_prime_1_27
-- reg_a = o1_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001011000000000100000000000000100001100110111",
--  (1473) square_with_reduction_special_prime_1_28
-- reg_a = a2_X; reg_b = a2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001011000000000100000000000000100001001000011",
--  (1474) square_with_reduction_special_prime_1_29
-- reg_a = o2_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
"000000100001011000000000100000000000000100001001010111",
--  (1475) square_with_reduction_special_prime_1_30
-- reg_a = o3_X; reg_b = primeSP1; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
"000000100001011000010000100000000000000100000101110111",
--  (1476) square_with_reduction_special_prime_1_31
-- reg_a = a2_X; reg_b = a3_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001011000000100100000100001000100001101000011",
--  (1477) square_with_reduction_special_prime_1_32
-- reg_a = o2_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001011000000000100000000000000100001101010111",
--  (1478) square_with_reduction_special_prime_1_33
-- reg_a = o3_X; reg_b = primeSP2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
"000000100001011000010000100000000000001000101001110111",
--  (1479) square_with_reduction_special_prime_1_34
-- reg_a = a3_X; reg_b = a3_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001011000000000100000100001100100001101100011",
--  (1480) square_with_reduction_special_prime_1_35
-- reg_a = o3_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; o3_X = reg_o >> 256; operation : a*b + acc;
"000000100001011001110000100000000000001101001101110111",
--  (1481) square_with_reduction_special_prime_1_36
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (1482) square_with_reduction_special_prime_1_37
-- -- In case of sizes 5, 6, 7, 8
-- reg_a = a0_X; reg_b = a3_X; reg_acc = reg_o; o3_X = reg_o; operation : 2*a*b + acc;
"000000100001100000010100100000000000010001101100000011",
--  (1483) square_with_reduction_special_prime_1_38
-- reg_a = o0_X; reg_b = primeSP4; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001100000000000100000100000000100010000010111",
--  (1484) square_with_reduction_special_prime_1_39
-- reg_a = a1_X; reg_b = a3_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001100000000100100000000000000100001100100011",
--  (1485) square_with_reduction_special_prime_1_40
-- reg_a = o1_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001100110111",
--  (1486) square_with_reduction_special_prime_1_41
-- reg_a = a2_X; reg_b = a2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001001000011",
--  (1487) square_with_reduction_special_prime_1_42
-- reg_a = o2_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001001010111",
--  (1488) square_with_reduction_special_prime_1_43
-- reg_a = o3_X; reg_b = primeSP1; reg_acc = reg_o; operation : a*b + acc;
"001001100001100000000000100000000000000100000101110111",
--  (1489) square_with_reduction_special_prime_1_44
-- -- In case of size 5
-- reg_a = a0_X; reg_b = a4_X; reg_acc = reg_o; o4_X = reg_o; Enable sign b; operation : 2*a*b + acc;
"000000100001100000010100100000000001010110010000000011",
--  (1490) square_with_reduction_special_prime_1_45
-- reg_a = a1_X; reg_b = a4_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001100000000100100000100001000100010000100011",
--  (1491) square_with_reduction_special_prime_1_46
-- reg_a = o1_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100010000110111",
--  (1492) square_with_reduction_special_prime_1_47
-- reg_a = a2_X; reg_b = a3_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001100000000100100000000000000100001101000011",
--  (1493) square_with_reduction_special_prime_1_48
-- reg_a = o2_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001101010111",
--  (1494) square_with_reduction_special_prime_1_49
-- reg_a = o3_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001001110111",
--  (1495) square_with_reduction_special_prime_1_50
-- reg_a = o4_X; reg_b = primeSP1; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
"000000100001100000010000100000000000000100000110010111",
--  (1496) square_with_reduction_special_prime_1_51
-- reg_a = a2_X; reg_b = a4_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001100000000100100000100001000100010001000011",
--  (1497) square_with_reduction_special_prime_1_52
-- reg_a = o2_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100010001010111",
--  (1498) square_with_reduction_special_prime_1_53
-- reg_a = a3_X; reg_b = a3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001101100011",
--  (1499) square_with_reduction_special_prime_1_54
-- reg_a = o3_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001101110111",
--  (1500) square_with_reduction_special_prime_1_55
-- reg_a = o4_X; reg_b = primeSP2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
"000000100001100000010000100000000000001000101010010111",
--  (1501) square_with_reduction_special_prime_1_56
-- reg_a = a3_X; reg_b = a4_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001100000000100100000100001000100010001100011",
--  (1502) square_with_reduction_special_prime_1_57
-- reg_a = o3_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100010001110111",
--  (1503) square_with_reduction_special_prime_1_58
-- reg_a = o4_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
"000000100001100000010000100000000000001101001110010111",
--  (1504) square_with_reduction_special_prime_1_59
-- reg_a = a4_X; reg_b = a4_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001100000000000100000100001100100010010000011",
--  (1505) square_with_reduction_special_prime_1_60
-- reg_a = o4_X; reg_b = primeSP4; reg_acc = reg_o; o3_X = reg_o; o4_X = reg_o >> 256; operation : a*b + acc;
"000000100001100001110000100000000000010001110010010111",
--  (1506) square_with_reduction_special_prime_1_61
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (1507) square_with_reduction_special_prime_1_62
-- -- In case of sizes 6, 7, 8
-- reg_a = a0_X; reg_b = a4_X; reg_acc = reg_o; o4_X = reg_o; operation : 2*a*b + acc;
"000000100001101000010100100000000000010110010000000011",
--  (1508) square_with_reduction_special_prime_1_63
-- reg_a = o0_X; reg_b = primeSP5; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001101000000000100000100000000100010100010111",
--  (1509) square_with_reduction_special_prime_1_64
-- reg_a = a1_X; reg_b = a4_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001101000000100100000000000000100010000100011",
--  (1510) square_with_reduction_special_prime_1_65
-- reg_a = o1_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010000110111",
--  (1511) square_with_reduction_special_prime_1_66
-- reg_a = a2_X; reg_b = a3_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001101000000100100000000000000100001101000011",
--  (1512) square_with_reduction_special_prime_1_67
-- reg_a = o2_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001101010111",
--  (1513) square_with_reduction_special_prime_1_68
-- reg_a = o3_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001001110111",
--  (1514) square_with_reduction_special_prime_1_69
-- reg_a = o4_X; reg_b = primeSP1; reg_acc = reg_o; operation : a*b + acc;
"001101100001101000000000100000000000000100000110010111",
--  (1515) square_with_reduction_special_prime_1_70
-- -- In case of size 6
-- reg_a = a0_X; reg_b = a5_X; reg_acc = reg_o; o5_X = reg_o; Enable sign b; operation : 2*a*b + acc;
"000000100001101000010100100000000001010010110100000011",
--  (1516) square_with_reduction_special_prime_1_71
-- reg_a = a1_X; reg_b = a5_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001101000000100100000100001000100010100100011",
--  (1517) square_with_reduction_special_prime_1_72
-- reg_a = o1_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010100110111",
--  (1518) square_with_reduction_special_prime_1_73
-- reg_a = a2_X; reg_b = a4_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001101000000100100000000000000100010001000011",
--  (1519) square_with_reduction_special_prime_1_74
-- reg_a = o2_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010001010111",
--  (1520) square_with_reduction_special_prime_1_75
-- reg_a = a3_X; reg_b = a3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001101100011",
--  (1521) square_with_reduction_special_prime_1_76
-- reg_a = o3_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001101110111",
--  (1522) square_with_reduction_special_prime_1_77
-- reg_a = o4_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001010010111",
--  (1523) square_with_reduction_special_prime_1_78
-- reg_a = o5_X; reg_b = primeSP1; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
"000000100001101000010000100000000000000100000110110111",
--  (1524) square_with_reduction_special_prime_1_79
-- reg_a = a2_X; reg_b = a5_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001101000000100100000100001000100010101000011",
--  (1525) square_with_reduction_special_prime_1_80
-- reg_a = o2_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010101010111",
--  (1526) square_with_reduction_special_prime_1_81
-- reg_a = a3_X; reg_b = a4_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001101000000100100000000000000100010001100011",
--  (1527) square_with_reduction_special_prime_1_82
-- reg_a = o3_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010001110111",
--  (1528) square_with_reduction_special_prime_1_83
-- reg_a = o4_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001110010111",
--  (1529) square_with_reduction_special_prime_1_84
-- reg_a = o5_X; reg_b = primeSP2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
"000000100001101000010000100000000000001000101010110111",
--  (1530) square_with_reduction_special_prime_1_85
-- reg_a = a3_X; reg_b = a5_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001101000000100100000100001000100010101100011",
--  (1531) square_with_reduction_special_prime_1_86
-- reg_a = o3_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010101110111",
--  (1532) square_with_reduction_special_prime_1_87
-- reg_a = a4_X; reg_b = a4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010010000011",
--  (1533) square_with_reduction_special_prime_1_88
-- reg_a = o4_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010010010111",
--  (1534) square_with_reduction_special_prime_1_89
-- reg_a = o5_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
"000000100001101000010000100000000000001101001110110111",
--  (1535) square_with_reduction_special_prime_1_90
-- reg_a = a4_X; reg_b = a5_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001101000000100100000100001000100010110000011",
--  (1536) square_with_reduction_special_prime_1_91
-- reg_a = o4_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010110010111",
--  (1537) square_with_reduction_special_prime_1_92
-- reg_a = o5_X; reg_b = primeSP4; reg_acc = reg_o; o3_X = reg_o; operation : a*b + acc;
"000000100001101000010000100000000000010001110010110111",
--  (1538) square_with_reduction_special_prime_1_93
-- reg_a = a5_X; reg_b = a5_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001101000000000100000100001100100010110100011",
--  (1539) square_with_reduction_special_prime_1_94
-- reg_a = o5_X; reg_b = primeSP5; reg_acc = reg_o; o4_X = reg_o; o5_X = reg_o >> 256; operation : a*b + acc;
"000000100001101001110000100000000000010110010110110111",
--  (1540) square_with_reduction_special_prime_1_95
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (1541) square_with_reduction_special_prime_1_96
-- -- In case of sizes 7, 8
-- reg_a = a0_X; reg_b = a5_X; reg_acc = reg_o; o5_X = reg_o; operation : 2*a*b + acc;
"000000100001110000010100100000000000011010110100000011",
--  (1542) square_with_reduction_special_prime_1_97
-- reg_a = o0_X; reg_b = primeSP6; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001110000000000100000100000000100011000010111",
--  (1543) square_with_reduction_special_prime_1_98
-- reg_a = a1_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001110000000100100000000000000100010100100011",
--  (1544) square_with_reduction_special_prime_1_99
-- reg_a = o1_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010100110111",
--  (1545) square_with_reduction_special_prime_1_100
-- reg_a = a2_X; reg_b = a4_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001110000000100100000000000000100010001000011",
--  (1546) square_with_reduction_special_prime_1_101
-- reg_a = o2_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010001010111",
--  (1547) square_with_reduction_special_prime_1_102
-- reg_a = a3_X; reg_b = a3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001101100011",
--  (1548) square_with_reduction_special_prime_1_103
-- reg_a = o3_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001101110111",
--  (1549) square_with_reduction_special_prime_1_104
-- reg_a = o4_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001010010111",
--  (1550) square_with_reduction_special_prime_1_105
-- reg_a = o5_X; reg_b = primeSP1; reg_acc = reg_o; operation : a*b + acc;
"010010000001110000000000100000000000000100000110110111",
--  (1551) square_with_reduction_special_prime_1_106
-- -- In case of size 7
-- reg_a = a0_X; reg_b = a6_X; reg_acc = reg_o; o6_X = reg_o; Enable sign b; operation : 2*a*b + acc;
"000000100001110000010100100000000001011111011000000011",
--  (1552) square_with_reduction_special_prime_1_107
-- reg_a = a1_X; reg_b = a6_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001110000000100100000100001000100011000100011",
--  (1553) square_with_reduction_special_prime_1_108
-- reg_a = o1_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100011000110111",
--  (1554) square_with_reduction_special_prime_1_109
-- reg_a = a2_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001110000000100100000000000000100010101000011",
--  (1555) square_with_reduction_special_prime_1_110
-- reg_a = o2_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010101010111",
--  (1556) square_with_reduction_special_prime_1_111
-- reg_a = a3_X; reg_b = a4_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001110000000100100000000000000100010001100011",
--  (1557) square_with_reduction_special_prime_1_112
-- reg_a = o3_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010001110111",
--  (1558) square_with_reduction_special_prime_1_113
-- reg_a = o4_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001110010111",
--  (1559) square_with_reduction_special_prime_1_114
-- reg_a = o5_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001010110111",
--  (1560) square_with_reduction_special_prime_1_115
-- reg_a = o6_X; reg_b = primeSP1; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
"000000100001110000010000100000000000000100000111010111",
--  (1561) square_with_reduction_special_prime_1_116
-- reg_a = a2_X; reg_b = a6_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001110000000100100000100001000100011001000011",
--  (1562) square_with_reduction_special_prime_1_117
-- reg_a = o2_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100011001010111",
--  (1563) square_with_reduction_special_prime_1_118
-- reg_a = a3_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001110000000100100000000000000100010101100011",
--  (1564) square_with_reduction_special_prime_1_119
-- reg_a = o3_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010101110111",
--  (1565) square_with_reduction_special_prime_1_120
-- reg_a = a4_X; reg_b = a4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010010000011",
--  (1566) square_with_reduction_special_prime_1_121
-- reg_a = o4_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010010010111",
--  (1567) square_with_reduction_special_prime_1_122
-- reg_a = o5_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001110110111",
--  (1568) square_with_reduction_special_prime_1_123
-- reg_a = o6_X; reg_b = primeSP2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
"000000100001110000010000100000000000001000101011010111",
--  (1569) square_with_reduction_special_prime_1_124
-- reg_a = a3_X; reg_b = a6_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001110000000100100000100001000100011001100011",
--  (1570) square_with_reduction_special_prime_1_125
-- reg_a = o3_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100011001110111",
--  (1571) square_with_reduction_special_prime_1_126
-- reg_a = a4_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001110000000100100000000000000100010110000011",
--  (1572) square_with_reduction_special_prime_1_127
-- reg_a = o4_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010110010111",
--  (1573) square_with_reduction_special_prime_1_128
-- reg_a = o5_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010010110111",
--  (1574) square_with_reduction_special_prime_1_129
-- reg_a = o6_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
"000000100001110000010000100000000000001101001111010111",
--  (1575) square_with_reduction_special_prime_1_130
-- reg_a = a4_X; reg_b = a6_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001110000000100100000100001000100011010000011",
--  (1576) square_with_reduction_special_prime_1_131
-- reg_a = o4_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100011010010111",
--  (1577) square_with_reduction_special_prime_1_132
-- reg_a = a5_X; reg_b = a5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010110100011",
--  (1578) square_with_reduction_special_prime_1_133
-- reg_a = o5_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010110110111",
--  (1579) square_with_reduction_special_prime_1_134
-- reg_a = o6_X; reg_b = primeSP4; reg_acc = reg_o; o3_X = reg_o; operation : a*b + acc;
"000000100001110000010000100000000000010001110011010111",
--  (1580) square_with_reduction_special_prime_1_135
-- reg_a = a5_X; reg_b = a6_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001110000000100100000100001000100011010100011",
--  (1581) square_with_reduction_special_prime_1_136
-- reg_a = o5_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100011010110111",
--  (1582) square_with_reduction_special_prime_1_137
-- reg_a = o6_X; reg_b = primeSP5; reg_acc = reg_o; o4_X = reg_o; operation : a*b + acc;
"000000100001110000010000100000000000010110010111010111",
--  (1583) square_with_reduction_special_prime_1_138
-- reg_a = a6_X; reg_b = a6_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001110000000000100000100001100100011011000011",
--  (1584) square_with_reduction_special_prime_1_139
-- reg_a = o6_X; reg_b = primeSP6; reg_acc = reg_o; o5_X = reg_o; o6_X = reg_o >> 256; operation : a*b + acc;
"000000100001110001110000100000000000011010111011010111",
--  (1585) square_with_reduction_special_prime_1_140
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (1586) square_with_reduction_special_prime_1_141
-- -- In case of size 8
-- reg_a = a0_X; reg_b = a6_X; reg_acc = reg_o; o6_X = reg_o; operation : 2*a*b + acc;
"000000100001111000010100100000000000011111011000000011",
--  (1587) square_with_reduction_special_prime_1_142
-- reg_a = o0_X; reg_b = primeSP7; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001111000000000100000100000000100011100010111",
--  (1588) square_with_reduction_special_prime_1_143
-- reg_a = a1_X; reg_b = a6_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001111000000100100000000000000100011000100011",
--  (1589) square_with_reduction_special_prime_1_144
-- reg_a = o1_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011000110111",
--  (1590) square_with_reduction_special_prime_1_145
-- reg_a = a2_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001111000000100100000000000000100010101000011",
--  (1591) square_with_reduction_special_prime_1_146
-- reg_a = o2_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010101010111",
--  (1592) square_with_reduction_special_prime_1_147
-- reg_a = a3_X; reg_b = a4_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001111000000100100000000000000100010001100011",
--  (1593) square_with_reduction_special_prime_1_148
-- reg_a = o3_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010001110111",
--  (1594) square_with_reduction_special_prime_1_149
-- reg_a = o4_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001110010111",
--  (1595) square_with_reduction_special_prime_1_150
-- reg_a = o5_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001010110111",
--  (1596) square_with_reduction_special_prime_1_151
-- reg_a = o6_X; reg_b = primeSP1; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100000111010111",
--  (1597) square_with_reduction_special_prime_1_152
-- reg_a = a0_X; reg_b = a7_X; reg_acc = reg_o; o7_X = reg_o; Enable sign b; operation : 2*a*b + acc;
"000000100001111000010100100000000001000011111100000011",
--  (1598) square_with_reduction_special_prime_1_153
-- reg_a = a1_X; reg_b = a7_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001111000000100100000100001000100011100100011",
--  (1599) square_with_reduction_special_prime_1_154
-- reg_a = o1_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011100110111",
--  (1600) square_with_reduction_special_prime_1_155
-- reg_a = a2_X; reg_b = a6_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001111000000100100000000000000100011001000011",
--  (1601) square_with_reduction_special_prime_1_156
-- reg_a = o2_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011001010111",
--  (1602) square_with_reduction_special_prime_1_157
-- reg_a = a3_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001111000000100100000000000000100010101100011",
--  (1603) square_with_reduction_special_prime_1_158
-- reg_a = o3_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010101110111",
--  (1604) square_with_reduction_special_prime_1_159
-- reg_a = a4_X; reg_b = a4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010010000011",
--  (1605) square_with_reduction_special_prime_1_160
-- reg_a = o4_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010010010111",
--  (1606) square_with_reduction_special_prime_1_161
-- reg_a = o5_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001110110111",
--  (1607) square_with_reduction_special_prime_1_162
-- reg_a = o6_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001011010111",
--  (1608) square_with_reduction_special_prime_1_163
-- reg_a = o7_X; reg_b = primeSP1; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000000100000111110111",
--  (1609) square_with_reduction_special_prime_1_164
-- reg_a = a2_X; reg_b = a7_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001111000000100100000100001000100011101000011",
--  (1610) square_with_reduction_special_prime_1_165
-- reg_a = o2_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011101010111",
--  (1611) square_with_reduction_special_prime_1_166
-- reg_a = a3_X; reg_b = a6_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001111000000100100000000000000100011001100011",
--  (1612) square_with_reduction_special_prime_1_167
-- reg_a = o3_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011001110111",
--  (1613) square_with_reduction_special_prime_1_168
-- reg_a = a4_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001111000000100100000000000000100010110000011",
--  (1614) square_with_reduction_special_prime_1_169
-- reg_a = o4_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010110010111",
--  (1615) square_with_reduction_special_prime_1_170
-- reg_a = o5_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010010110111",
--  (1616) square_with_reduction_special_prime_1_171
-- reg_a = o6_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001111010111",
--  (1617) square_with_reduction_special_prime_1_172
-- reg_a = o7_X; reg_b = primeSP2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000001000101011110111",
--  (1618) square_with_reduction_special_prime_1_173
-- reg_a = a3_X; reg_b = a7_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001111000000100100000100001000100011101100011",
--  (1619) square_with_reduction_special_prime_1_174
-- reg_a = o3_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011101110111",
--  (1620) square_with_reduction_special_prime_1_175
-- reg_a = a4_X; reg_b = a6_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001111000000100100000000000000100011010000011",
--  (1621) square_with_reduction_special_prime_1_176
-- reg_a = o4_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011010010111",
--  (1622) square_with_reduction_special_prime_1_177
-- reg_a = a5_X; reg_b = a5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010110100011",
--  (1623) square_with_reduction_special_prime_1_178
-- reg_a = o5_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010110110111",
--  (1624) square_with_reduction_special_prime_1_179
-- reg_a = o6_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010011010111",
--  (1625) square_with_reduction_special_prime_1_180
-- reg_a = o7_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000001101001111110111",
--  (1626) square_with_reduction_special_prime_1_181
-- reg_a = a4_X; reg_b = a7_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001111000000100100000100001000100011110000011",
--  (1627) square_with_reduction_special_prime_1_182
-- reg_a = o4_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011110010111",
--  (1628) square_with_reduction_special_prime_1_183
-- reg_a = a5_X; reg_b = a6_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001111000000100100000000000000100011010100011",
--  (1629) square_with_reduction_special_prime_1_184
-- reg_a = o5_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011010110111",
--  (1630) square_with_reduction_special_prime_1_185
-- reg_a = o6_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010111010111",
--  (1631) square_with_reduction_special_prime_1_186
-- reg_a = o7_X; reg_b = primeSP4; reg_acc = reg_o; o3_X = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000010001110011110111",
--  (1632) square_with_reduction_special_prime_1_187
-- reg_a = a5_X; reg_b = a7_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001111000000100100000100001000100011110100011",
--  (1633) square_with_reduction_special_prime_1_188
-- reg_a = o5_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011110110111",
--  (1634) square_with_reduction_special_prime_1_189
-- reg_a = a6_X; reg_b = a6_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011011000011",
--  (1635) square_with_reduction_special_prime_1_190
-- reg_a = o6_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011011010111",
--  (1636) square_with_reduction_special_prime_1_191
-- reg_a = o7_X; reg_b = primeSP5; reg_acc = reg_o; o4_X = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000010110010111110111",
--  (1637) square_with_reduction_special_prime_1_192
-- reg_a = a6_X; reg_b = a7_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001111000000100100000100001000100011111000011",
--  (1638) square_with_reduction_special_prime_1_193
-- reg_a = o6_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011111010111",
--  (1639) square_with_reduction_special_prime_1_194
-- reg_a = o7_X; reg_b = primeSP6; reg_acc = reg_o; o5_X = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000011010111011110111",
--  (1640) square_with_reduction_special_prime_1_195
-- reg_a = a7_X; reg_b = a7_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001111000000000100000100001100100011111100011",
--  (1641) square_with_reduction_special_prime_1_196
-- reg_a = o7_X; reg_b = primeSP7; reg_acc = reg_o; o6_X = reg_o; o7_X = reg_o >> 256; operation : a*b + acc;
"000000100001111001110000100000000000011111011111110111",
--  (1642) square_with_reduction_special_prime_1_197
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (1643) square_with_reduction_special_prime_2_0
-- -- In case of size 2, 3, 4, 5, 6, 7, 8
-- reg_a = a0_X; reg_b = a0_X; reg_acc = 0; o0_X = reg_o; operation : a*b + acc;
"000010000001001000010000100000010000000100000000000011",
--  (1644) square_with_reduction_special_prime_2_1
-- -- In case of size 2
-- reg_a = a0_X; reg_b = a1_X; reg_acc = reg_o; o1_X = reg_o; Enable sign b; operation : 2*a*b + acc;
"000000100001001000010100100000000001001000100100000011",
--  (1645) square_with_reduction_special_prime_2_2
-- reg_a = a1_X; reg_b = a1_X; reg_acc = reg_o >> 256; Enable sign a,b; o0_X = reg_o; o1_X = reg_o >> 256; operation : a*b + acc;
"000000100001001001110000100000100001100100000100100011",
--  (1646) square_with_reduction_special_prime_2_3
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (1647) square_with_reduction_special_prime_2_4
-- -- In case of size 3, 4, 5, 6, 7, 8
-- reg_a = a0_X; reg_b = a1_X; reg_acc = reg_o >> 256; o1_X = reg_o; operation : 2*a*b + acc;
"000000100001010000010100100000100000001000100100000011",
--  (1648) square_with_reduction_special_prime_2_5
-- reg_a = o0_X; reg_b = primeSP2; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001010000000000100000100000000100001000010111",
--  (1649) square_with_reduction_special_prime_2_6
-- reg_a = a1_X; reg_b = a1_X; reg_acc = reg_o; operation : a*b + acc;
"000011100001010000000000100000000000000100000100100011",
--  (1650) square_with_reduction_special_prime_2_7
-- -- In case of size 3
-- reg_a = a0_X; reg_b = a2_X; reg_acc = reg_o; o2_X = reg_o; Enable sign b; operation : 2*a*b + acc;
"000000100001010000010100100000000001001101001000000011",
--  (1651) square_with_reduction_special_prime_2_8
-- reg_a = a1_X; reg_b = a2_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001010000000100100000100001000100001000100011",
--  (1652) square_with_reduction_special_prime_2_9
-- reg_a = o1_X; reg_b = primeSP2; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
"000000100001010000010000100000000000000100001000110111",
--  (1653) square_with_reduction_special_prime_2_10
-- reg_a = a2_X; reg_b = a2_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001010000000000100000100001100100001001000011",
--  (1654) square_with_reduction_special_prime_2_11
-- reg_a = o2_X; reg_b = primeSP2; reg_acc = reg_o; o1_X = reg_o; o2_X = reg_o >> 256; operation : a*b + acc;
"000000100001010001110000100000000000001000101001010111",
--  (1655) square_with_reduction_special_prime_2_12
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (1656) square_with_reduction_special_prime_2_13
-- -- In case of size 4, 5, 6, 7, 8
-- reg_a = a0_X; reg_b = a2_X; reg_acc = reg_o; o2_X = reg_o; operation : 2*a*b + acc;
"000000100001011000010100100000000000001101001000000011",
--  (1657) square_with_reduction_special_prime_2_14
-- reg_a = o0_X; reg_b = primeSP3; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001011000000000100000100000000100001100010111",
--  (1658) square_with_reduction_special_prime_2_15
-- reg_a = a1_X; reg_b = a2_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001011000000100100000000000000100001000100011",
--  (1659) square_with_reduction_special_prime_2_16
-- reg_a = o1_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
"000110000001011000000000100000000000000100001000110111",
--  (1660) square_with_reduction_special_prime_2_17
-- -- In case of size 4
-- reg_a = a0_X; reg_b = a3_X; reg_acc = reg_o; o3_X = reg_o; Enable sign b; operation : 2*a*b + acc;
"000000100001011000010100100000000001010001101100000011",
--  (1661) square_with_reduction_special_prime_2_18
-- reg_a = a1_X; reg_b = a3_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001011000000100100000100001000100001100100011",
--  (1662) square_with_reduction_special_prime_2_19
-- reg_a = o1_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001011000000000100000000000000100001100110111",
--  (1663) square_with_reduction_special_prime_2_20
-- reg_a = a2_X; reg_b = a2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001011000000000100000000000000100001001000011",
--  (1664) square_with_reduction_special_prime_2_21
-- reg_a = o2_X; reg_b = primeSP2; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
"000000100001011000010000100000000000000100001001010111",
--  (1665) square_with_reduction_special_prime_2_22
-- reg_a = a2_X; reg_b = a3_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001011000000100100000100001000100001101000011",
--  (1666) square_with_reduction_special_prime_2_23
-- reg_a = o2_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001011000000000100000000000000100001101010111",
--  (1667) square_with_reduction_special_prime_2_24
-- reg_a = o3_X; reg_b = primeSP2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
"000000100001011000010000100000000000001000101001110111",
--  (1668) square_with_reduction_special_prime_2_25
-- reg_a = a3_X; reg_b = a3_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001011000000000100000100001100100001101100011",
--  (1669) square_with_reduction_special_prime_2_26
-- reg_a = o3_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; o3_X = reg_o >> 256; operation : a*b + acc;
"000000100001011001110000100000000000001101001101110111",
--  (1670) square_with_reduction_special_prime_2_27
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (1671) square_with_reduction_special_prime_2_28
-- -- In case of size 5, 6, 7, 8
-- reg_a = a0_X; reg_b = a3_X; reg_acc = reg_o; o3_X = reg_o; operation : 2*a*b + acc;
"000000100001100000010100100000000000010001101100000011",
--  (1672) square_with_reduction_special_prime_2_29
-- reg_a = o0_X; reg_b = primeSP4; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001100000000000100000100000000100010000010111",
--  (1673) square_with_reduction_special_prime_2_30
-- reg_a = a1_X; reg_b = a3_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001100000000100100000000000000100001100100011",
--  (1674) square_with_reduction_special_prime_2_31
-- reg_a = o1_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001100110111",
--  (1675) square_with_reduction_special_prime_2_32
-- reg_a = a2_X; reg_b = a2_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001001000011",
--  (1676) square_with_reduction_special_prime_2_33
-- reg_a = o2_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
"001001000001100000000000100000000000000100001001010111",
--  (1677) square_with_reduction_special_prime_2_34
-- -- In case of size 5
-- reg_a = a0_X; reg_b = a4_X; reg_acc = reg_o; o4_X = reg_o; Enable sign b; operation : 2*a*b + acc;
"000000100001100000010100100000000001010110010000000011",
--  (1678) square_with_reduction_special_prime_2_35
-- reg_a = a1_X; reg_b = a4_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001100000000100100000100001000100010000100011",
--  (1679) square_with_reduction_special_prime_2_36
-- reg_a = o1_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100010000110111",
--  (1680) square_with_reduction_special_prime_2_37
-- reg_a = a2_X; reg_b = a3_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001100000000100100000000000000100001101000011",
--  (1681) square_with_reduction_special_prime_2_38
-- reg_a = o2_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001101010111",
--  (1682) square_with_reduction_special_prime_2_39
-- reg_a = o3_X; reg_b = primeSP2; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
"000000100001100000010000100000000000000100001001110111",
--  (1683) square_with_reduction_special_prime_2_40
-- reg_a = a2_X; reg_b = a4_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001100000000100100000100001000100010001000011",
--  (1684) square_with_reduction_special_prime_2_41
-- reg_a = o2_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100010001010111",
--  (1685) square_with_reduction_special_prime_2_42
-- reg_a = a3_X; reg_b = a3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001101100011",
--  (1686) square_with_reduction_special_prime_2_43
-- reg_a = o3_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001101110111",
--  (1687) square_with_reduction_special_prime_2_44
-- reg_a = o4_X; reg_b = primeSP2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
"000000100001100000010000100000000000001000101010010111",
--  (1688) square_with_reduction_special_prime_2_45
-- reg_a = a3_X; reg_b = a4_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001100000000100100000100001000100010001100011",
--  (1689) square_with_reduction_special_prime_2_46
-- reg_a = o3_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100010001110111",
--  (1690) square_with_reduction_special_prime_2_47
-- reg_a = o4_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
"000000100001100000010000100000000000001101001110010111",
--  (1691) square_with_reduction_special_prime_2_48
-- reg_a = a4_X; reg_b = a4_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001100000000000100000100001100100010010000011",
--  (1692) square_with_reduction_special_prime_2_49
-- reg_a = o4_X; reg_b = primeSP4; reg_acc = reg_o; o3_X = reg_o; o4_X = reg_o >> 256; operation : a*b + acc;
"000000100001100001110000100000000000010001110010010111",
--  (1693) square_with_reduction_special_prime_2_50
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (1694) square_with_reduction_special_prime_2_51
-- -- In case of sizes 6, 7, 8
-- reg_a = a0_X; reg_b = a4_X; reg_acc = reg_o; o4_X = reg_o; operation : 2*a*b + acc;
"000000100001101000010100100000000000010110010000000011",
--  (1695) square_with_reduction_special_prime_2_52
-- reg_a = o0_X; reg_b = primeSP5; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001101000000000100000100000000100010100010111",
--  (1696) square_with_reduction_special_prime_2_53
-- reg_a = a1_X; reg_b = a4_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001101000000100100000000000000100010000100011",
--  (1697) square_with_reduction_special_prime_2_54
-- reg_a = o1_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010000110111",
--  (1698) square_with_reduction_special_prime_2_55
-- reg_a = a2_X; reg_b = a3_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001101000000100100000000000000100001101000011",
--  (1699) square_with_reduction_special_prime_2_56
-- reg_a = o2_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001101010111",
--  (1700) square_with_reduction_special_prime_2_57
-- reg_a = o3_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
"001101000001101000000000100000000000000100001001110111",
--  (1701) square_with_reduction_special_prime_2_58
-- -- In case of size 6
-- reg_a = a0_X; reg_b = a5_X; reg_acc = reg_o; o5_X = reg_o; Enable sign b; operation : 2*a*b + acc;
"000000100001101000010100100000000001011010110100000011",
--  (1702) square_with_reduction_special_prime_2_59
-- reg_a = a1_X; reg_b = a5_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001101000000100100000100001000100010100100011",
--  (1703) square_with_reduction_special_prime_2_60
-- reg_a = o1_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010100110111",
--  (1704) square_with_reduction_special_prime_2_61
-- reg_a = a2_X; reg_b = a4_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001101000000100100000000000000100010001000011",
--  (1705) square_with_reduction_special_prime_2_62
-- reg_a = o2_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010001010111",
--  (1706) square_with_reduction_special_prime_2_63
-- reg_a = a3_X; reg_b = a3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001101100011",
--  (1707) square_with_reduction_special_prime_2_64
-- reg_a = o3_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001101110111",
--  (1708) square_with_reduction_special_prime_2_65
-- reg_a = o4_X; reg_b = primeSP2; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
"000000100001101000010000100000000000000100001010010111",
--  (1709) square_with_reduction_special_prime_2_66
-- reg_a = a2_X; reg_b = a5_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001101000000100100000100001000100010101000011",
--  (1710) square_with_reduction_special_prime_2_67
-- reg_a = o2_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010101010111",
--  (1711) square_with_reduction_special_prime_2_68
-- reg_a = a3_X; reg_b = a4_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001101000000100100000000000000100010001100011",
--  (1712) square_with_reduction_special_prime_2_69
-- reg_a = o3_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010001110111",
--  (1713) square_with_reduction_special_prime_2_70
-- reg_a = o4_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001110010111",
--  (1714) square_with_reduction_special_prime_2_71
-- reg_a = o5_X; reg_b = primeSP2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
"000000100001101000010000100000000000001000101010110111",
--  (1715) square_with_reduction_special_prime_2_72
-- reg_a = a3_X; reg_b = a5_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001101000000100100000100001000100010101100011",
--  (1716) square_with_reduction_special_prime_2_73
-- reg_a = o3_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010101110111",
--  (1717) square_with_reduction_special_prime_2_74
-- reg_a = a4_X; reg_b = a4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010010000011",
--  (1718) square_with_reduction_special_prime_2_75
-- reg_a = o4_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010010010111",
--  (1719) square_with_reduction_special_prime_2_76
-- reg_a = o5_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
"000000100001101000010000100000000000001101001110110111",
--  (1720) square_with_reduction_special_prime_2_77
-- reg_a = a4_X; reg_b = a5_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001101000000100100000100001000100010110000011",
--  (1721) square_with_reduction_special_prime_2_78
-- reg_a = o4_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010110010111",
--  (1722) square_with_reduction_special_prime_2_79
-- reg_a = o5_X; reg_b = primeSP4; reg_acc = reg_o; o3_X = reg_o; operation : a*b + acc;
"000000100001101000010000100000000000010001110010110111",
--  (1723) square_with_reduction_special_prime_2_80
-- reg_a = a5_X; reg_b = a5_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001101000000000100000100001100100010110100011",
--  (1724) square_with_reduction_special_prime_2_81
-- reg_a = o5_X; reg_b = primeSP5; reg_acc = reg_o; o4_X = reg_o; o5_X = reg_o >> 256; operation : a*b + acc;
"000000100001101001110000100000000000010110010110110111",
--  (1725) square_with_reduction_special_prime_2_82
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (1726) square_with_reduction_special_prime_2_83
-- -- In case of sizes 7, 8
-- reg_a = a0_X; reg_b = a5_X; reg_acc = reg_o; o5_X = reg_o; operation : 2*a*b + acc;
"000000100001110000010100100000000000011010110100000011",
--  (1727) square_with_reduction_special_prime_2_84
-- reg_a = o0_X; reg_b = primeSP6; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001110000000000100000100000000100011000010111",
--  (1728) square_with_reduction_special_prime_2_85
-- reg_a = a1_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001110000000100100000000000000100010100100011",
--  (1729) square_with_reduction_special_prime_2_86
-- reg_a = o1_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010100110111",
--  (1730) square_with_reduction_special_prime_2_87
-- reg_a = a2_X; reg_b = a4_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001110000000100100000000000000100010001000011",
--  (1731) square_with_reduction_special_prime_2_88
-- reg_a = o2_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010001010111",
--  (1732) square_with_reduction_special_prime_2_89
-- reg_a = a3_X; reg_b = a3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001101100011",
--  (1733) square_with_reduction_special_prime_2_90
-- reg_a = o3_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001101110111",
--  (1734) square_with_reduction_special_prime_2_91
-- reg_a = o4_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
"010001100001110000000000100000000000000100001010010111",
--  (1735) square_with_reduction_special_prime_2_92
-- -- In case of size 7
-- reg_a = a0_X; reg_b = a6_X; reg_acc = reg_o; o6_X = reg_o; Enable sign b; operation : 2*a*b + acc;
"000000100001110000010100100000000001011111011000000011",
--  (1736) square_with_reduction_special_prime_2_93
-- reg_a = a1_X; reg_b = a6_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001110000000100100000100001000100011000100011",
--  (1737) square_with_reduction_special_prime_2_94
-- reg_a = o1_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100011000110111",
--  (1738) square_with_reduction_special_prime_2_95
-- reg_a = a2_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001110000000100100000000000000100010101000011",
--  (1739) square_with_reduction_special_prime_2_96
-- reg_a = o2_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010101010111",
--  (1740) square_with_reduction_special_prime_2_97
-- reg_a = a3_X; reg_b = a4_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001110000000100100000000000000100010001100011",
--  (1741) square_with_reduction_special_prime_2_98
-- reg_a = o3_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010001110111",
--  (1742) square_with_reduction_special_prime_2_99
-- reg_a = o4_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001110010111",
--  (1743) square_with_reduction_special_prime_2_100
-- reg_a = o5_X; reg_b = primeSP2; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
"000000100001110000010000100000000000000100001010110111",
--  (1744) square_with_reduction_special_prime_2_101
-- reg_a = a2_X; reg_b = a6_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001110000000100100000100001000100011001000011",
--  (1745) square_with_reduction_special_prime_2_102
-- reg_a = o2_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100011001010111",
--  (1746) square_with_reduction_special_prime_2_103
-- reg_a = a3_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001110000000100100000000000000100010101100011",
--  (1747) square_with_reduction_special_prime_2_104
-- reg_a = o3_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010101110111",
--  (1748) square_with_reduction_special_prime_2_105
-- reg_a = a4_X; reg_b = a4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010010000011",
--  (1749) square_with_reduction_special_prime_2_106
-- reg_a = o4_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010010010111",
--  (1750) square_with_reduction_special_prime_2_107
-- reg_a = o5_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001110110111",
--  (1751) square_with_reduction_special_prime_2_108
-- reg_a = o6_X; reg_b = primeSP2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
"000000100001110000010000100000000000001000101011010111",
--  (1752) square_with_reduction_special_prime_2_109
-- reg_a = a3_X; reg_b = a6_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001110000000100100000100001000100011001100011",
--  (1753) square_with_reduction_special_prime_2_110
-- reg_a = o3_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100011001110111",
--  (1754) square_with_reduction_special_prime_2_111
-- reg_a = a4_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001110000000100100000000000000100010110000011",
--  (1755) square_with_reduction_special_prime_2_112
-- reg_a = o4_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010110010111",
--  (1756) square_with_reduction_special_prime_2_113
-- reg_a = o5_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010010110111",
--  (1757) square_with_reduction_special_prime_2_114
-- reg_a = o6_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
"000000100001110000010000100000000000001101001111010111",
--  (1758) square_with_reduction_special_prime_2_115
-- reg_a = a4_X; reg_b = a6_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001110000000100100000100001000100011010000011",
--  (1759) square_with_reduction_special_prime_2_116
-- reg_a = o4_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100011010010111",
--  (1760) square_with_reduction_special_prime_2_117
-- reg_a = a5_X; reg_b = a5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010110100011",
--  (1761) square_with_reduction_special_prime_2_118
-- reg_a = o5_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010110110111",
--  (1762) square_with_reduction_special_prime_2_119
-- reg_a = o6_X; reg_b = primeSP4; reg_acc = reg_o; o3_X = reg_o; operation : a*b + acc;
"000000100001110000010000100000000000010001110011010111",
--  (1763) square_with_reduction_special_prime_2_120
-- reg_a = a5_X; reg_b = a6_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001110000000100100000100001000100011010100011",
--  (1764) square_with_reduction_special_prime_2_121
-- reg_a = o5_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100011010110111",
--  (1765) square_with_reduction_special_prime_2_122
-- reg_a = o6_X; reg_b = primeSP5; reg_acc = reg_o; o4_X = reg_o; operation : a*b + acc;
"000000100001110000010000100000000000010110010111010111",
--  (1766) square_with_reduction_special_prime_2_123
-- reg_a = a6_X; reg_b = a6_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001110000000000100000100001100100011011000011",
--  (1767) square_with_reduction_special_prime_2_124
-- reg_a = o6_X; reg_b = primeSP6; reg_acc = reg_o; o5_X = reg_o; o6_X = reg_o >> 256; operation : a*b + acc;
"000000100001110001110000100000000000011010111011010111",
--  (1768) square_with_reduction_special_prime_2_125
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (1769) square_with_reduction_special_prime_2_126
-- -- In case of size 8
-- reg_a = a0_X; reg_b = a6_X; reg_acc = reg_o; o6_X = reg_o; operation : 2*a*b + acc;
"000000100001111000010100100000000000011111011000000011",
--  (1770) square_with_reduction_special_prime_2_127
-- reg_a = o0_X; reg_b = primeSP7; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001111000000000100000100000000100011100010111",
--  (1771) square_with_reduction_special_prime_2_128
-- reg_a = a1_X; reg_b = a6_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001111000000100100000000000000100011000100011",
--  (1772) square_with_reduction_special_prime_2_129
-- reg_a = o1_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011000110111",
--  (1773) square_with_reduction_special_prime_2_130
-- reg_a = a2_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001111000000100100000000000000100010101000011",
--  (1774) square_with_reduction_special_prime_2_131
-- reg_a = o2_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010101010111",
--  (1775) square_with_reduction_special_prime_2_132
-- reg_a = a3_X; reg_b = a4_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001111000000100100000000000000100010001100011",
--  (1776) square_with_reduction_special_prime_2_133
-- reg_a = o3_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010001110111",
--  (1777) square_with_reduction_special_prime_2_134
-- reg_a = o4_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001110010111",
--  (1778) square_with_reduction_special_prime_2_135
-- reg_a = o5_X; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001010110111",
--  (1779) square_with_reduction_special_prime_2_136
-- reg_a = a0_X; reg_b = a7_X; reg_acc = reg_o; o7_X = reg_o; Enable sign b; operation : 2*a*b + acc;
"000000100001111000010100100000000001000011111100000011",
--  (1780) square_with_reduction_special_prime_2_137
-- reg_a = a1_X; reg_b = a7_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001111000000100100000100001000100011100100011",
--  (1781) square_with_reduction_special_prime_2_138
-- reg_a = o1_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011100110111",
--  (1782) square_with_reduction_special_prime_2_139
-- reg_a = a2_X; reg_b = a6_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001111000000100100000000000000100011001000011",
--  (1783) square_with_reduction_special_prime_2_140
-- reg_a = o2_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011001010111",
--  (1784) square_with_reduction_special_prime_2_141
-- reg_a = a3_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001111000000100100000000000000100010101100011",
--  (1785) square_with_reduction_special_prime_2_142
-- reg_a = o3_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010101110111",
--  (1786) square_with_reduction_special_prime_2_143
-- reg_a = a4_X; reg_b = a4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010010000011",
--  (1787) square_with_reduction_special_prime_2_144
-- reg_a = o4_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010010010111",
--  (1788) square_with_reduction_special_prime_2_145
-- reg_a = o5_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001110110111",
--  (1789) square_with_reduction_special_prime_2_146
-- reg_a = o6_X; reg_b = primeSP2; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000000100001011010111",
--  (1790) square_with_reduction_special_prime_2_147
-- reg_a = a2_X; reg_b = a7_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001111000000100100000100001000100011101000011",
--  (1791) square_with_reduction_special_prime_2_148
-- reg_a = o2_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011101010111",
--  (1792) square_with_reduction_special_prime_2_149
-- reg_a = a3_X; reg_b = a6_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001111000000100100000000000000100011001100011",
--  (1793) square_with_reduction_special_prime_2_150
-- reg_a = o3_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011001110111",
--  (1794) square_with_reduction_special_prime_2_151
-- reg_a = a4_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001111000000100100000000000000100010110000011",
--  (1795) square_with_reduction_special_prime_2_152
-- reg_a = o4_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010110010111",
--  (1796) square_with_reduction_special_prime_2_153
-- reg_a = o5_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010010110111",
--  (1797) square_with_reduction_special_prime_2_154
-- reg_a = o6_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001111010111",
--  (1798) square_with_reduction_special_prime_2_155
-- reg_a = o7_X; reg_b = primeSP2; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000001000101011110111",
--  (1799) square_with_reduction_special_prime_2_156
-- reg_a = a3_X; reg_b = a7_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001111000000100100000100001000100011101100011",
--  (1800) square_with_reduction_special_prime_2_157
-- reg_a = o3_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011101110111",
--  (1801) square_with_reduction_special_prime_2_158
-- reg_a = a4_X; reg_b = a6_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001111000000100100000000000000100011010000011",
--  (1802) square_with_reduction_special_prime_2_159
-- reg_a = o4_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011010010111",
--  (1803) square_with_reduction_special_prime_2_160
-- reg_a = a5_X; reg_b = a5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010110100011",
--  (1804) square_with_reduction_special_prime_2_161
-- reg_a = o5_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010110110111",
--  (1805) square_with_reduction_special_prime_2_162
-- reg_a = o6_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010011010111",
--  (1806) square_with_reduction_special_prime_2_163
-- reg_a = o7_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000001101001111110111",
--  (1807) square_with_reduction_special_prime_2_164
-- reg_a = a4_X; reg_b = a7_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001111000000100100000100001000100011110000011",
--  (1808) square_with_reduction_special_prime_2_165
-- reg_a = o4_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011110010111",
--  (1809) square_with_reduction_special_prime_2_166
-- reg_a = a5_X; reg_b = a6_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001111000000100100000000000000100011010100011",
--  (1810) square_with_reduction_special_prime_2_167
-- reg_a = o5_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011010110111",
--  (1811) square_with_reduction_special_prime_2_168
-- reg_a = o6_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010111010111",
--  (1812) square_with_reduction_special_prime_2_169
-- reg_a = o7_X; reg_b = primeSP4; reg_acc = reg_o; o3_X = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000010001110011110111",
--  (1813) square_with_reduction_special_prime_2_170
-- reg_a = a5_X; reg_b = a7_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001111000000100100000100001000100011110100011",
--  (1814) square_with_reduction_special_prime_2_171
-- reg_a = o5_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011110110111",
--  (1815) square_with_reduction_special_prime_2_172
-- reg_a = a6_X; reg_b = a6_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011011000011",
--  (1816) square_with_reduction_special_prime_2_173
-- reg_a = o6_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011011010111",
--  (1817) square_with_reduction_special_prime_2_174
-- reg_a = o7_X; reg_b = primeSP5; reg_acc = reg_o; o4_X = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000010110010111110111",
--  (1818) square_with_reduction_special_prime_2_175
-- reg_a = a6_X; reg_b = a7_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001111000000100100000100001000100011111000011",
--  (1819) square_with_reduction_special_prime_2_176
-- reg_a = o6_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011111010111",
--  (1820) square_with_reduction_special_prime_2_177
-- reg_a = o7_X; reg_b = primeSP6; reg_acc = reg_o; o5_X = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000011010111011110111",
--  (1821) square_with_reduction_special_prime_2_178
-- reg_a = a7_X; reg_b = a7_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001111000000000100000100001100100011111100011",
--  (1822) square_with_reduction_special_prime_2_179
-- reg_a = o7_X; reg_b = primeSP7; reg_acc = reg_o; o6_X = reg_o; o7_X = reg_o >> 256; operation : a*b + acc;
"000000100001111001110000100000000000011111011111110111",
--  (1823) square_with_reduction_special_prime_2_180
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (1824) square_with_reduction_special_prime_3_0
-- -- In case of sizes 3, 4, 5, 6, 7, 8
-- reg_a = a0_X; reg_b = a0_X; reg_acc = 0; o0_X = reg_o; operation : a*b + acc;
"000000100001010000010000100000010000000100000000000011",
--  (1825) square_with_reduction_special_prime_3_1
-- reg_a = a0_X; reg_b = a1_X; reg_acc = reg_o >> 256; o1_X = reg_o; operation : 2*a*b + acc;
"000000100001010000010100100000100000001000100100000011",
--  (1826) square_with_reduction_special_prime_3_2
-- reg_a = a1_X; reg_b = a1_X; reg_acc = reg_o >> 256; operation : a*b + acc;
"000010100001010000000000100000100000000100000100100011",
--  (1827) square_with_reduction_special_prime_3_3
-- -- In case of size 3
-- reg_a = a0_X; reg_b = a2_X; reg_acc = reg_o; o2_X = reg_o; Enable sign b; operation : 2*a*b + acc;
"000000100001010000010100100000000001001101001000000011",
--  (1828) square_with_reduction_special_prime_3_4
-- reg_a = a1_X; reg_b = a2_X; reg_acc = reg_o >> 256; Enable sign b; o0_X = reg_o; operation : 2*a*b + acc;
"000000100001010000010100100000100001000100001000100011",
--  (1829) square_with_reduction_special_prime_3_5
-- reg_a = a2_X; reg_b = a2_X; reg_acc = reg_o >> 256; Enable sign a,b; o1_X = reg_o; o2_X = reg_o >> 256; operation : a*b + acc;
"000000100001010001110000100000100001101000101001000011",
--  (1830) square_with_reduction_special_prime_3_6
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (1831) square_with_reduction_special_prime_3_7
-- -- In case of sizes 4, 5, 6, 7, 8
-- reg_a = a0_X; reg_b = a2_X; reg_acc = reg_o; o2_X = reg_o; operation : 2*a*b + acc;
"000000100001011000010100100000000000001101001000000011",
--  (1832) square_with_reduction_special_prime_3_8
-- reg_a = o0_X; reg_b = primeSP3; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001011000000000100000100000000100001100010111",
--  (1833) square_with_reduction_special_prime_3_9
-- reg_a = a1_X; reg_b = a2_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000101000001011000000100100000000000000100001000100011",
--  (1834) square_with_reduction_special_prime_3_10
-- -- In case of size 4
-- reg_a = a0_X; reg_b = a3_X; reg_acc = reg_o; o3_X = reg_o; Enable sign b; operation : 2*a*b + acc;
"000000100001011000010100100000000001010001101100000011",
--  (1835) square_with_reduction_special_prime_3_11
-- reg_a = a1_X; reg_b = a3_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001011000000100100000100001000100001100100011",
--  (1836) square_with_reduction_special_prime_3_12
-- reg_a = o1_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001011000000000100000000000000100001100110111",
--  (1837) square_with_reduction_special_prime_3_13
-- reg_a = a2_X; reg_b = a2_X; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
"000000100001011000010000100000000000000100001001000011",
--  (1838) square_with_reduction_special_prime_3_14
-- reg_a = a2_X; reg_b = a3_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001011000000100100000100001000100001101000011",
--  (1839) square_with_reduction_special_prime_3_15
-- reg_a = o2_X; reg_b = primeSP3; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
"000000100001011000010000100000000000001000101101010111",
--  (1840) square_with_reduction_special_prime_3_16
-- reg_a = a3_X; reg_b = a3_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001011000000000100000100001100100001101100011",
--  (1841) square_with_reduction_special_prime_3_17
-- reg_a = o3_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; o3_X = reg_o >> 256; operation : a*b + acc;
"000000100001011001110000100000000000001101001101110111",
--  (1842) square_with_reduction_special_prime_3_18
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (1843) square_with_reduction_special_prime_3_19
-- -- In case of sizes 5, 6, 7, 8
-- reg_a = a0_X; reg_b = a3_X; reg_acc = reg_o; o3_X = reg_o; operation : 2*a*b + acc;
"000000100001100000010100100000000000010001101100000011",
--  (1844) square_with_reduction_special_prime_3_20
-- reg_a = o0_X; reg_b = primeSP4; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001100000000000100000100000000100010000010111",
--  (1845) square_with_reduction_special_prime_3_21
-- reg_a = a1_X; reg_b = a3_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001100000000100100000000000000100001100100011",
--  (1846) square_with_reduction_special_prime_3_22
-- reg_a = o1_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001100110111",
--  (1847) square_with_reduction_special_prime_3_23
-- reg_a = a2_X; reg_b = a2_X; reg_acc = reg_o; operation : a*b + acc;
"001000000001100000000000100000000000000100001001000011",
--  (1848) square_with_reduction_special_prime_3_24
-- -- In case of size 5
-- reg_a = a0_X; reg_b = a4_X; reg_acc = reg_o; o4_X = reg_o; Enable sign b; operation : 2*a*b + acc;
"000000100001100000010100100000000001010110010000000011",
--  (1849) square_with_reduction_special_prime_3_25
-- reg_a = a1_X; reg_b = a4_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001100000000100100000100001000100010000100011",
--  (1850) square_with_reduction_special_prime_3_26
-- reg_a = o1_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100010000110111",
--  (1851) square_with_reduction_special_prime_3_27
-- reg_a = a2_X; reg_b = a3_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001100000000100100000000000000100001101000011",
--  (1852) square_with_reduction_special_prime_3_28
-- reg_a = o2_X; reg_b = primeSP3; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
"000000100001100000010000100000000000000100001101010111",
--  (1853) square_with_reduction_special_prime_3_29
-- reg_a = a2_X; reg_b = a4_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001100000000100100000100001000100010001000011",
--  (1854) square_with_reduction_special_prime_3_30
-- reg_a = o2_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100010001010111",
--  (1855) square_with_reduction_special_prime_3_31
-- reg_a = a3_X; reg_b = a3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100001101100011",
--  (1856) square_with_reduction_special_prime_3_32
-- reg_a = o3_X; reg_b = primeSP3; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
"000000100001100000010000100000000000001000101101110111",
--  (1857) square_with_reduction_special_prime_3_33
-- reg_a = a3_X; reg_b = a4_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001100000000100100000100001000100010001100011",
--  (1858) square_with_reduction_special_prime_3_34
-- reg_a = o3_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001100000000000100000000000000100010001110111",
--  (1859) square_with_reduction_special_prime_3_35
-- reg_a = o4_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
"000000100001100000010000100000000000001101001110010111",
--  (1860) square_with_reduction_special_prime_3_36
-- reg_a = a4_X; reg_b = a4_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001100000000000100000100001100100010010000011",
--  (1861) square_with_reduction_special_prime_3_37
-- reg_a = o4_X; reg_b = primeSP4; reg_acc = reg_o; o3_X = reg_o; o4_X = reg_o >> 256; operation : a*b + acc;
"000000100001100001110000100000000000010001110010010111",
--  (1862) square_with_reduction_special_prime_3_38
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (1863) square_with_reduction_special_prime_3_39
-- -- In case of sizes 6, 7, 8
-- reg_a = a0_X; reg_b = a4_X; reg_acc = reg_o; o4_X = reg_o; operation : 2*a*b + acc;
"000000100001101000010100100000000000010110010000000011",
--  (1864) square_with_reduction_special_prime_3_40
-- reg_a = o0_X; reg_b = primeSP5; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001101000000000100000100000000100010100010111",
--  (1865) square_with_reduction_special_prime_3_41
-- reg_a = a1_X; reg_b = a4_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001101000000100100000000000000100010000100011",
--  (1866) square_with_reduction_special_prime_3_42
-- reg_a = o1_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010000110111",
--  (1867) square_with_reduction_special_prime_3_43
-- reg_a = a2_X; reg_b = a3_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001101000000100100000000000000100001101000011",
--  (1868) square_with_reduction_special_prime_3_44
-- reg_a = o2_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"001100000001101000000000100000000000000100001101010111",
--  (1869) square_with_reduction_special_prime_3_45
-- -- In case of size 6
-- reg_a = a0_X; reg_b = a5_X; reg_acc = reg_o; o5_X = reg_o; Enable sign b; operation : 2*a*b + acc;
"000000100001101000010100100000000001011010110100000011",
--  (1870) square_with_reduction_special_prime_3_46
-- reg_a = a1_X; reg_b = a5_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001101000000100100000100001000100010100100011",
--  (1871) square_with_reduction_special_prime_3_47
-- reg_a = o1_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010100110111",
--  (1872) square_with_reduction_special_prime_3_48
-- reg_a = a2_X; reg_b = a4_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001101000000100100000000000000100010001000011",
--  (1873) square_with_reduction_special_prime_3_49
-- reg_a = o2_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010001010111",
--  (1874) square_with_reduction_special_prime_3_50
-- reg_a = a3_X; reg_b = a3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100001101100011",
--  (1875) square_with_reduction_special_prime_3_51
-- reg_a = o3_X; reg_b = primeSP3; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
"000000100001101000010000100000000000000100001101110111",
--  (1876) square_with_reduction_special_prime_3_52
-- reg_a = a2_X; reg_b = a5_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001101000000100100000100001000100010101000011",
--  (1877) square_with_reduction_special_prime_3_53
-- reg_a = o2_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010101010111",
--  (1878) square_with_reduction_special_prime_3_54
-- reg_a = a3_X; reg_b = a4_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001101000000100100000000000000100010001100011",
--  (1879) square_with_reduction_special_prime_3_55
-- reg_a = o3_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010001110111",
--  (1880) square_with_reduction_special_prime_3_56
-- reg_a = o4_X; reg_b = primeSP3; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
"000000100001101000010000100000000000001000101110010111",
--  (1881) square_with_reduction_special_prime_3_57
-- reg_a = a3_X; reg_b = a5_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001101000000100100000100001000100010101100011",
--  (1882) square_with_reduction_special_prime_3_58
-- reg_a = o3_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010101110111",
--  (1883) square_with_reduction_special_prime_3_59
-- reg_a = a4_X; reg_b = a4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010010000011",
--  (1884) square_with_reduction_special_prime_3_60
-- reg_a = o4_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010010010111",
--  (1885) square_with_reduction_special_prime_3_61
-- reg_a = o5_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
"000000100001101000010000100000000000001101001110110111",
--  (1886) square_with_reduction_special_prime_3_62
-- reg_a = a4_X; reg_b = a5_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001101000000100100000100001000100010110000011",
--  (1887) square_with_reduction_special_prime_3_63
-- reg_a = o4_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001101000000000100000000000000100010110010111",
--  (1888) square_with_reduction_special_prime_3_64
-- reg_a = o5_X; reg_b = primeSP4; reg_acc = reg_o; o3_X = reg_o; operation : a*b + acc;
"000000100001101000010000100000000000010001110010110111",
--  (1889) square_with_reduction_special_prime_3_65
-- reg_a = a5_X; reg_b = a5_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001101000000000100000100001100100010110100011",
--  (1890) square_with_reduction_special_prime_3_66
-- reg_a = o5_X; reg_b = primeSP5; reg_acc = reg_o; o4_X = reg_o; o5_X = reg_o >> 256; operation : a*b + acc;
"000000100001101001110000100000000000010110010110110111",
--  (1891) square_with_reduction_special_prime_3_67
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (1892) square_with_reduction_special_prime_3_68
-- -- In case of sizes 7, 8
-- reg_a = a0_X; reg_b = a5_X; reg_acc = reg_o; o5_X = reg_o; operation : 2*a*b + acc;
"000000100001110000010100100000000000011010110100000011",
--  (1893) square_with_reduction_special_prime_3_69
-- reg_a = o0_X; reg_b = primeSP6; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001110000000000100000100000000100011000010111",
--  (1894) square_with_reduction_special_prime_3_70
-- reg_a = a1_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001110000000100100000000000000100010100100011",
--  (1895) square_with_reduction_special_prime_3_71
-- reg_a = o1_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010100110111",
--  (1896) square_with_reduction_special_prime_3_72
-- reg_a = a2_X; reg_b = a4_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001110000000100100000000000000100010001000011",
--  (1897) square_with_reduction_special_prime_3_73
-- reg_a = o2_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010001010111",
--  (1898) square_with_reduction_special_prime_3_74
-- reg_a = a3_X; reg_b = a3_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100001101100011",
--  (1899) square_with_reduction_special_prime_3_75
-- reg_a = o3_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"010000100001110000000000100000000000000100001101110111",
--  (1900) square_with_reduction_special_prime_3_76
-- -- In case of size 7
-- reg_a = a0_X; reg_b = a6_X; reg_acc = reg_o; o6_X = reg_o; Enable sign b; operation : 2*a*b + acc;
"000000100001110000010100100000000001011111011000000011",
--  (1901) square_with_reduction_special_prime_3_77
-- reg_a = a1_X; reg_b = a6_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001110000000100100000100001000100011000100011",
--  (1902) square_with_reduction_special_prime_3_78
-- reg_a = o1_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100011000110111",
--  (1903) square_with_reduction_special_prime_3_79
-- reg_a = a2_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001110000000100100000000000000100010101000011",
--  (1904) square_with_reduction_special_prime_3_80
-- reg_a = o2_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010101010111",
--  (1905) square_with_reduction_special_prime_3_81
-- reg_a = a3_X; reg_b = a4_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001110000000100100000000000000100010001100011",
--  (1906) square_with_reduction_special_prime_3_82
-- reg_a = o3_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010001110111",
--  (1907) square_with_reduction_special_prime_3_83
-- reg_a = o4_X; reg_b = primeSP3; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
"000000100001110000010000100000000000000100001110010111",
--  (1908) square_with_reduction_special_prime_3_84
-- reg_a = a2_X; reg_b = a6_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001110000000100100000100001000100011001000011",
--  (1909) square_with_reduction_special_prime_3_85
-- reg_a = o2_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100011001010111",
--  (1910) square_with_reduction_special_prime_3_86
-- reg_a = a3_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001110000000100100000000000000100010101100011",
--  (1911) square_with_reduction_special_prime_3_87
-- reg_a = o3_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010101110111",
--  (1912) square_with_reduction_special_prime_3_88
-- reg_a = a4_X; reg_b = a4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010010000011",
--  (1913) square_with_reduction_special_prime_3_89
-- reg_a = o4_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010010010111",
--  (1914) square_with_reduction_special_prime_3_90
-- reg_a = o5_X; reg_b = primeSP3; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
"000000100001110000010000100000000000001000101110110111",
--  (1915) square_with_reduction_special_prime_3_91
-- reg_a = a3_X; reg_b = a6_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001110000000100100000100001000100011001100011",
--  (1916) square_with_reduction_special_prime_3_92
-- reg_a = o3_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100011001110111",
--  (1917) square_with_reduction_special_prime_3_93
-- reg_a = a4_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001110000000100100000000000000100010110000011",
--  (1918) square_with_reduction_special_prime_3_94
-- reg_a = o4_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010110010111",
--  (1919) square_with_reduction_special_prime_3_95
-- reg_a = o5_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010010110111",
--  (1920) square_with_reduction_special_prime_3_96
-- reg_a = o6_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
"000000100001110000010000100000000000001101001111010111",
--  (1921) square_with_reduction_special_prime_3_97
-- reg_a = a4_X; reg_b = a6_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001110000000100100000100001000100011010000011",
--  (1922) square_with_reduction_special_prime_3_98
-- reg_a = o4_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100011010010111",
--  (1923) square_with_reduction_special_prime_3_99
-- reg_a = a5_X; reg_b = a5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010110100011",
--  (1924) square_with_reduction_special_prime_3_100
-- reg_a = o5_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100010110110111",
--  (1925) square_with_reduction_special_prime_3_101
-- reg_a = o6_X; reg_b = primeSP4; reg_acc = reg_o; o3_X = reg_o; operation : a*b + acc;
"000000100001110000010000100000000000010001110011010111",
--  (1926) square_with_reduction_special_prime_3_102
-- reg_a = a5_X; reg_b = a6_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001110000000100100000100001000100011010100011",
--  (1927) square_with_reduction_special_prime_3_103
-- reg_a = o5_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001110000000000100000000000000100011010110111",
--  (1928) square_with_reduction_special_prime_3_104
-- reg_a = o6_X; reg_b = primeSP5; reg_acc = reg_o; o4_X = reg_o; operation : a*b + acc;
"000000100001110000010000100000000000010110010111010111",
--  (1929) square_with_reduction_special_prime_3_105
-- reg_a = a6_X; reg_b = a6_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001110000000000100000100001100100011011000011",
--  (1930) square_with_reduction_special_prime_3_106
-- reg_a = o6_X; reg_b = primeSP6; reg_acc = reg_o; o5_X = reg_o; o6_X = reg_o >> 256; operation : a*b + acc;
"000000100001110001110000100000000000011010111011010111",
--  (1931) square_with_reduction_special_prime_3_107
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (1932) square_with_reduction_special_prime_3_108
-- -- In case of size 8
-- reg_a = a0_X; reg_b = a6_X; reg_acc = reg_o; o6_X = reg_o; operation : 2*a*b + acc;
"000000100001111000010100100000000000011011011000000011",
--  (1933) square_with_reduction_special_prime_3_109
-- reg_a = o0_X; reg_b = primeSP7; reg_acc = reg_o >> 256; operation : a*b + acc;
"000000100001111000000000100000100000000100011100010111",
--  (1934) square_with_reduction_special_prime_3_110
-- reg_a = a1_X; reg_b = a6_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001111000000100100000000000000100011000100011",
--  (1935) square_with_reduction_special_prime_3_111
-- reg_a = o1_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011000110111",
--  (1936) square_with_reduction_special_prime_3_112
-- reg_a = a2_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001111000000100100000000000000100010101000011",
--  (1937) square_with_reduction_special_prime_3_113
-- reg_a = o2_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010101010111",
--  (1938) square_with_reduction_special_prime_3_114
-- reg_a = a3_X; reg_b = a4_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001111000000100100000000000000100010001100011",
--  (1939) square_with_reduction_special_prime_3_115
-- reg_a = o3_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010001110111",
--  (1940) square_with_reduction_special_prime_3_116
-- reg_a = o4_X; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100001110010111",
--  (1941) square_with_reduction_special_prime_3_117
-- reg_a = a0_X; reg_b = a7_X; reg_acc = reg_o; o7_X = reg_o; Enable sign b; operation : 2*a*b + acc;
"000000100001111000010100100000000001011111111100000011",
--  (1942) square_with_reduction_special_prime_3_118
-- reg_a = a1_X; reg_b = a7_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001111000000100100000100001000100011100100011",
--  (1943) square_with_reduction_special_prime_3_119
-- reg_a = o1_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011100110111",
--  (1944) square_with_reduction_special_prime_3_120
-- reg_a = a2_X; reg_b = a6_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001111000000100100000000000000100011001000011",
--  (1945) square_with_reduction_special_prime_3_121
-- reg_a = o2_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011001010111",
--  (1946) square_with_reduction_special_prime_3_122
-- reg_a = a3_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001111000000100100000000000000100010101100011",
--  (1947) square_with_reduction_special_prime_3_123
-- reg_a = o3_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010101110111",
--  (1948) square_with_reduction_special_prime_3_124
-- reg_a = a4_X; reg_b = a4_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010010000011",
--  (1949) square_with_reduction_special_prime_3_125
-- reg_a = o4_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010010010111",
--  (1950) square_with_reduction_special_prime_3_126
-- reg_a = o5_X; reg_b = primeSP3; reg_acc = reg_o; o0_X = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000000100001110110111",
--  (1951) square_with_reduction_special_prime_3_127
-- reg_a = a2_X; reg_b = a7_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001111000000100100000100001000100011101000011",
--  (1952) square_with_reduction_special_prime_3_128
-- reg_a = o2_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011101010111",
--  (1953) square_with_reduction_special_prime_3_129
-- reg_a = a3_X; reg_b = a6_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001111000000100100000000000000100011001100011",
--  (1954) square_with_reduction_special_prime_3_130
-- reg_a = o3_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011001110111",
--  (1955) square_with_reduction_special_prime_3_131
-- reg_a = a4_X; reg_b = a5_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001111000000100100000000000000100010110000011",
--  (1956) square_with_reduction_special_prime_3_132
-- reg_a = o4_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010110010111",
--  (1957) square_with_reduction_special_prime_3_133
-- reg_a = o5_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010010110111",
--  (1958) square_with_reduction_special_prime_3_134
-- reg_a = o6_X; reg_b = primeSP3; reg_acc = reg_o; o1_X = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000001000101111010111",
--  (1959) square_with_reduction_special_prime_3_135
-- reg_a = a3_X; reg_b = a7_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001111000000100100000100001000100011101100011",
--  (1960) square_with_reduction_special_prime_3_136
-- reg_a = o3_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011101110111",
--  (1961) square_with_reduction_special_prime_3_137
-- reg_a = a4_X; reg_b = a6_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001111000000100100000000000000100011010000011",
--  (1962) square_with_reduction_special_prime_3_138
-- reg_a = o4_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011010010111",
--  (1963) square_with_reduction_special_prime_3_139
-- reg_a = a5_X; reg_b = a5_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010110100011",
--  (1964) square_with_reduction_special_prime_3_140
-- reg_a = o5_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010110110111",
--  (1965) square_with_reduction_special_prime_3_141
-- reg_a = o6_X; reg_b = primeSP4; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010011010111",
--  (1966) square_with_reduction_special_prime_3_142
-- reg_a = o7_X; reg_b = primeSP3; reg_acc = reg_o; o2_X = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000001101001111110111",
--  (1967) square_with_reduction_special_prime_3_143
-- reg_a = a4_X; reg_b = a7_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001111000000100100000100001000100011110000011",
--  (1968) square_with_reduction_special_prime_3_144
-- reg_a = o4_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011110010111",
--  (1969) square_with_reduction_special_prime_3_145
-- reg_a = a5_X; reg_b = a6_X; reg_acc = reg_o; operation : 2*a*b + acc;
"000000100001111000000100100000000000000100011010100011",
--  (1970) square_with_reduction_special_prime_3_146
-- reg_a = o5_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011010110111",
--  (1971) square_with_reduction_special_prime_3_147
-- reg_a = o6_X; reg_b = primeSP5; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100010111010111",
--  (1972) square_with_reduction_special_prime_3_148
-- reg_a = o7_X; reg_b = primeSP4; reg_acc = reg_o; o3_X = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000010001110011110111",
--  (1973) square_with_reduction_special_prime_3_149
-- reg_a = a5_X; reg_b = a7_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001111000000100100000100001000100011110100011",
--  (1974) square_with_reduction_special_prime_3_150
-- reg_a = o5_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011110110111",
--  (1975) square_with_reduction_special_prime_3_151
-- reg_a = a6_X; reg_b = a6_X; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011011000011",
--  (1976) square_with_reduction_special_prime_3_152
-- reg_a = o6_X; reg_b = primeSP6; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011011010111",
--  (1977) square_with_reduction_special_prime_3_153
-- reg_a = o7_X; reg_b = primeSP5; reg_acc = reg_o; o4_X = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000010110010111110111",
--  (1978) square_with_reduction_special_prime_3_154
-- reg_a = a6_X; reg_b = a7_X; reg_acc = reg_o >> 256; Enable sign b; operation : 2*a*b + acc;
"000000100001111000000100100000100001000100011111000011",
--  (1979) square_with_reduction_special_prime_3_155
-- reg_a = o6_X; reg_b = primeSP7; reg_acc = reg_o; operation : a*b + acc;
"000000100001111000000000100000000000000100011111010111",
--  (1980) square_with_reduction_special_prime_3_156
-- reg_a = o7_X; reg_b = primeSP6; reg_acc = reg_o; o5_X = reg_o; operation : a*b + acc;
"000000100001111000010000100000000000011010111011110111",
--  (1981) square_with_reduction_special_prime_3_157
-- reg_a = a7_X; reg_b = a7_X; reg_acc = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
"000000100001111000000000100000100001100100011111100011",
--  (1982) square_with_reduction_special_prime_3_158
-- reg_a = o7_X; reg_b = primeSP7; reg_acc = reg_o; o6_X = reg_o; o7_X = reg_o >> 256; operation : a*b + acc;
"000000100001111001110000100000000000011111011111110111",
--  (1983) square_with_reduction_special_prime_3_159
-- NOP 8 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
"000000000000000100000000100000011110000100000000000011",
--  (1984) addition_subtraction_direct_0
-- -- In case of size 1
-- reg_a = a0_X; reg_b = b0_X; reg_acc = 0; o0_0 = reg_o; Enable sign a,b; operation : b +/- a + acc;
"000000100001000000010000001000010001100100000000000010",
--  (1985) addition_subtraction_direct_1
-- NOP 4 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : b + a + acc;
"000000000000000100000000010000011110000100000000000010",
--  (1986) addition_subtraction_direct_2
-- -- In case of size 2, 3, 4, 5, 6, 7, 8
-- reg_a = a0_X; reg_b = b0_X; reg_acc = 0; o0_X = reg_o; operation : b +/- a + acc;
"000001100001001000010000001000010000000100000000000010",
--  (1987) addition_subtraction_direct_3
-- -- In case of size 2
-- reg_a = a1_X; reg_b = b1_X; reg_acc = reg_o >> 256; o1_X = reg_o; Enable sign a, b; operation : b +/- a + acc;
"000000100001001000010000001000100001101000100100100010",
--  (1988) addition_subtraction_direct_4
-- NOP 4 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : b + a + acc;
"000000000000000100000000010000011110000100000000000010",
--  (1989) addition_subtraction_direct_5
-- -- In case of size 3, 4, 5, 6, 7, 8
-- reg_a = a1_X; reg_b = b1_X; reg_acc = reg_o >> 256; o1_X = reg_o; operation : b +/- a + acc;
"000001100001010000010000001000100000001000100100100010",
--  (1990) addition_subtraction_direct_6
-- -- In case of size 3
-- reg_a = a2_X; reg_b = b2_X; reg_acc = reg_o >> 256; o2_X = reg_o; Enable sign a,b; operation : b +/- a + acc;
"000000100001010000010000001000100001100101001001000010",
--  (1991) addition_subtraction_direct_7
-- NOP 4 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : b + a + acc;
"000000000000000100000000010000011110000100000000000010",
--  (1992) addition_subtraction_direct_8
-- -- In case of size 4, 5, 6, 7, 8
-- reg_a = a2_X; reg_b = b2_X; reg_acc = reg_o >> 256; o2_X = reg_o; operation : b +/- a + acc;
"000001100001011000010000001000100000000101001001000010",
--  (1993) addition_subtraction_direct_9
-- -- In case of size 4
-- reg_a = a3_X; reg_b = b3_X; reg_acc = reg_o >> 256; o3_X = reg_o; Enable sign a,b; operation : b +/- a + acc;
"000000100001011000010000001000100001110001101101100010",
--  (1994) addition_subtraction_direct_10
-- NOP 4 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : b + a + acc;
"000000000000000100000000010000011110000100000000000010",
--  (1995) addition_subtraction_direct_11
-- -- In case of size 4, 5, 6, 7, 8
-- reg_a = a3_X; reg_b = b3_X; reg_acc = reg_o >> 256; o3_X = reg_o; operation : b +/- a + acc;
"000001100001100000010000001000100000010001101101100010",
--  (1996) addition_subtraction_direct_12
-- -- In case of size 5
-- reg_a = a4_X; reg_b = b4_X; reg_acc = reg_o >> 256; o4_X = reg_o; Enable sign a,b; operation : b +/- a + acc;
"000000100001100000010000001000100001110110010010000010",
--  (1997) addition_subtraction_direct_13
-- NOP 4 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : b + a + acc;
"000000000000000100000000010000011110000100000000000010",
--  (1998) addition_subtraction_direct_14
-- -- In case of size 6, 7, 8
-- reg_a = a4_X; reg_b = b4_X; reg_acc = reg_o >> 256; o4_X = reg_o; operation : b +/- a + acc;
"000001100001101000010000001000100000010110010010000010",
--  (1999) addition_subtraction_direct_15
-- -- In case of size 6
-- reg_a = a5_X; reg_b = b5_X; reg_acc = reg_o >> 256; o5_X = reg_o; Enable sign a,b; operation : b +/- a + acc;
"000000100001101000010000001000100001111010110110100010",
--  (2000) addition_subtraction_direct_16
-- NOP 4 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : b + a + acc;
"000000000000000100000000010000011110000100000000000010",
--  (2001) addition_subtraction_direct_17
-- -- In case of size 7, 8
-- reg_a = a5_X; reg_b = b5_X; reg_acc = reg_o >> 256; o5_X = reg_o; operation : b +/- a + acc;
"000001100001110000010000001000100000011010110110100010",
--  (2002) addition_subtraction_direct_18
-- -- In case of size 7
-- reg_a = a6_X; reg_b = b6_X; reg_acc = reg_o >> 256; o6_X = reg_o; Enable sign a,b; operation : b +/- a + acc;
"000000100001110000010000001000100001111111011011000010",
--  (2003) addition_subtraction_direct_19
-- NOP 4 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : b + a + acc;
"000000000000000100000000010000011110000100000000000010",
--  (2004) addition_subtraction_direct_20
-- -- In case of size 8
-- reg_a = a6_X; reg_b = b6_X; reg_acc = reg_o >> 256; o6_X = reg_o; operation : b +/- a + acc;
"000000100001111000010000001000100000011111011011000010",
--  (2005) addition_subtraction_direct_21
-- reg_a = a7_X; reg_b = b7_X; reg_acc = reg_o >> 256; o7_X = reg_o; Enable sign a,b; operation : b +/- a + acc;
"000000100001111000010000001000100001100011111111100010",
--  (2006) addition_subtraction_direct_22
-- NOP 4 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : b + a + acc;
"000000000000000100000000010000011110000100000000000010",
--  (2007) iterative_modular_reduction_0
-- -- In case of size 1
-- reg_a = a0_X; reg_b = 0; reg_acc = 0; Enable sign a,b; operation : b + a + acc;
"000000100001000000000000010000011001100100000000010010",
--  (2008) iterative_modular_reduction_1
-- reg_a = 0; reg_b = prime0; reg_acc = reg_o; reg_s = reg_o_positive; Enable sign a,b; operation : -s*b + a + acc
"000000100001000000000011000111000111100100000000010010",
--  (2009) iterative_modular_reduction_2
-- reg_a = 0; reg_b = prime0; reg_acc = reg_o; reg_s = reg_o_negative; Enable sign a,b; operation : s*b + a + acc
"000000100001000000000001010011000111100100000000010010",
--  (2010) iterative_modular_reduction_3
-- reg_a = 0; reg_b = prime0; reg_acc = reg_o; o0_X = reg_o; reg_s = reg_o_negative; Enable sign a,b; operation : s*b + a + acc
"000000100001000000010001010011000111100100000000010010",
--  (2011) iterative_modular_reduction_4
-- NOP 4 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : b + a + acc;
"000000000000000100000000010000011110000100000000000010",
--  (2012) iterative_modular_reduction_5
-- -- In case of size 2
-- reg_a = a1_X; reg_b = 0; reg_acc = 0; Enable sign a,b; operation : b + a + acc;
"000000100001001000000000010000011001100100000000110010",
--  (2013) iterative_modular_reduction_6
-- reg_a = a0_X; reg_b = prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_positive; operation : -s*b + a + acc
"000000100001001000010011000111010000000100000000010010",
--  (2014) iterative_modular_reduction_7
-- reg_a = a1_X; reg_b = prime1; reg_acc = reg_o >> 256; o1_X = reg_o; Enable sign a,b; operation : -s*b + a + acc
"000000100001001000010011000000100001101000100100110010",
--  (2015) iterative_modular_reduction_8
-- reg_a = o0_X; reg_b = prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc
"000000100001001000010001010011010000000100000000010110",
--  (2016) iterative_modular_reduction_9
-- reg_a = o1_X; reg_b = prime1; reg_acc = reg_o >> 256; o1_X = reg_o; Enable sign a,b operation : s*b + a + acc
"000000100001001000010001010000100001101000100100110110",
--  (2017) iterative_modular_reduction_10
-- reg_a = o0_X; reg_b = prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc
"000000100001001000010001010011010000000100000000010110",
--  (2018) iterative_modular_reduction_11
-- reg_a = o1_X; reg_b = prime1; reg_acc = reg_o >> 256; o1_X = reg_o; Enable sign a,b operation : s*b + a + acc
"000000100001001000010001010000100001101000100100110110",
--  (2019) iterative_modular_reduction_12
-- NOP 4 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : b + a + acc;
"000000000000000100000000010000011110000100000000000010",
--  (2020) iterative_modular_reduction_13
-- -- In case of size 3
-- reg_a = a2_X; reg_b = 0; reg_acc = 0; Enable sign a,b; operation : b + a + acc;
"000000100001010000000000010000011001101101001001010010",
--  (2021) iterative_modular_reduction_14
-- reg_a = a0_X; reg_b = prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_positive; operation : -s*b + a + acc
"000000100001010000010011000111010000000100000000010010",
--  (2022) iterative_modular_reduction_15
-- reg_a = a1_X; reg_b = prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : -s*b + a + acc
"000000100001010000010011000000100000001000100100110010",
--  (2023) iterative_modular_reduction_16
-- reg_a = a2_X; reg_b = prime2; reg_acc = reg_o >> 256; o2_X = reg_o; Enable sign a,b; operation : -s*b + a + acc
"000000100001010000010011000000100001101101001001010010",
--  (2024) iterative_modular_reduction_17
-- reg_a = o0_X; reg_b = prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc
"000000100001010000010001010011010000000100000000010110",
--  (2025) iterative_modular_reduction_18
-- reg_a = o1_X; reg_b = prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : s*b + a + acc
"000000100001010000010001010000100000001000100100110110",
--  (2026) iterative_modular_reduction_19
-- reg_a = o2_X; reg_b = prime2; reg_acc = reg_o >> 256; o2_X = reg_o; Enable sign a,b operation : s*b + a + acc
"000000100001010000010001010000100001101101001001010110",
--  (2027) iterative_modular_reduction_20
-- reg_a = o0_X; reg_b = prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc
"000000100001010000010001010011010000000100000000010110",
--  (2028) iterative_modular_reduction_21
-- reg_a = o1_X; reg_b = prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : s*b + a + acc
"000000100001010000010001010000100000001000100100110110",
--  (2029) iterative_modular_reduction_22
-- reg_a = o2_X; reg_b = prime2; reg_acc = reg_o >> 256; o2_X = reg_o; Enable sign a,b operation : s*b + a + acc
"000000100001010000010001010000100001101101001001010110",
--  (2030) iterative_modular_reduction_23
-- NOP 4 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : b + a + acc;
"000000000000000100000000010000011110000100000000000010",
--  (2031) iterative_modular_reduction_24
-- -- In case of size 4
-- reg_a = a3_X; reg_b = 0; reg_acc = 0; Enable sign a,b; operation : b + a + acc;
"000000100001011000000000010000011001100001101101110010",
--  (2032) iterative_modular_reduction_25
-- reg_a = a0_X; reg_b = prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_positive; operation : -s*b + a + acc
"000000100001011000010011000111010000000100000000010010",
--  (2033) iterative_modular_reduction_26
-- reg_a = a1_X; reg_b = prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : -s*b + a + acc
"000000100001011000010011000000100000001000100100110010",
--  (2034) iterative_modular_reduction_27
-- reg_a = a2_X; reg_b = prime2; reg_acc = reg_o >> 256; o2_X = reg_o; operation : -s*b + a + acc
"000000100001011000010011000000100000001101001001010010",
--  (2035) iterative_modular_reduction_28
-- reg_a = a3_X; reg_b = prime3; reg_acc = reg_o >> 256; o3_X = reg_o; Enable sign a,b; operation : -s*b + a + acc
"000000100001011000010011000000100001100001101101110010",
--  (2036) iterative_modular_reduction_29
-- reg_a = o0_X; reg_b = prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc
"000000100001011000010001010011010000000100000000010110",
--  (2037) iterative_modular_reduction_30
-- reg_a = o1_X; reg_b = prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : s*b + a + acc
"000000100001011000010001010000100000001000100100110110",
--  (2038) iterative_modular_reduction_31
-- reg_a = o2_X; reg_b = prime2; reg_acc = reg_o >> 256; o2_X = reg_o; operation : s*b + a + acc
"000000100001011000010001010000100000001101001001010110",
--  (2039) iterative_modular_reduction_32
-- reg_a = o3_X; reg_b = prime3; reg_acc = reg_o >> 256; o3_X = reg_o; Enable sign a,b; operation : s*b + a + acc
"000000100001011000010001010000100001100001101101110110",
--  (2040) iterative_modular_reduction_33
-- reg_a = o0_X; reg_b = prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc
"000000100001011000010001010011010000000100000000010110",
--  (2041) iterative_modular_reduction_34
-- reg_a = o1_X; reg_b = prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : s*b + a + acc
"000000100001011000010001010000100000001000100100110110",
--  (2042) iterative_modular_reduction_35
-- reg_a = o2_X; reg_b = prime2; reg_acc = reg_o >> 256; o2_X = reg_o; operation : s*b + a + acc
"000000100001011000010001010000100000001101001001010110",
--  (2043) iterative_modular_reduction_36
-- reg_a = o3_X; reg_b = prime3; reg_acc = reg_o >> 256; o3_X = reg_o; Enable sign a,b; operation : s*b + a + acc
"000000100001011000010001010000100001100001101101110110",
--  (2044) iterative_modular_reduction_37
-- NOP 4 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : b + a + acc;
"000000000000000100000000010000011110000100000000000010",
--  (2045) iterative_modular_reduction_38
-- -- In case of size 5
-- reg_a = a4_X; reg_b = 0; reg_acc = 0; Enable sign a,b; operation : b + a + acc;
"000000100001100000000000010000011001110110010010010010",
--  (2046) iterative_modular_reduction_39
-- reg_a = a0_X; reg_b = prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_positive; operation : -s*b + a + acc
"000000100001100000010011000111010000000100000000010010",
--  (2047) iterative_modular_reduction_40
-- reg_a = a1_X; reg_b = prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : -s*b + a + acc
"000000100001100000010011000000100000001000100100110010",
--  (2048) iterative_modular_reduction_41
-- reg_a = a2_X; reg_b = prime2; reg_acc = reg_o >> 256; o2_X = reg_o; operation : -s*b + a + acc
"000000100001100000010011000000100000001101001001010010",
--  (2049) iterative_modular_reduction_42
-- reg_a = a3_X; reg_b = prime3; reg_acc = reg_o >> 256; o3_X = reg_o; operation : -s*b + a + acc
"000000100001100000010011000000100000010001101101110010",
--  (2050) iterative_modular_reduction_43
-- reg_a = a4_X; reg_b = prime4; reg_acc = reg_o >> 256; o4_X = reg_o; Enable sign a,b; operation : -s*b + a + acc
"000000100001100000010011000000100001110110010010010010",
--  (2051) iterative_modular_reduction_44
-- reg_a = o0_X; reg_b = prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc
"000000100001100000010001010011010000000100000000010110",
--  (2052) iterative_modular_reduction_45
-- reg_a = o1_X; reg_b = prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : s*b + a + acc
"000000100001100000010001010000100000001000100100110110",
--  (2053) iterative_modular_reduction_46
-- reg_a = o2_X; reg_b = prime2; reg_acc = reg_o >> 256; o2_X = reg_o; operation : s*b + a + acc
"000000100001100000010001010000100000001101001001010110",
--  (2054) iterative_modular_reduction_47
-- reg_a = o3_X; reg_b = prime3; reg_acc = reg_o >> 256; o3_X = reg_o; operation : s*b + a + acc
"000000100001100000010001010000100000010001101101110110",
--  (2055) iterative_modular_reduction_48
-- reg_a = o4_X; reg_b = prime4; reg_acc = reg_o >> 256; o4_X = reg_o; Enable sign a,b; operation : s*b + a + acc
"000000100001100000010001010000100001110110010010010110",
--  (2056) iterative_modular_reduction_49
-- reg_a = o0_X; reg_b = prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc
"000000100001100000010001010011010000000100000000010110",
--  (2057) iterative_modular_reduction_50
-- reg_a = o1_X; reg_b = prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : s*b + a + acc
"000000100001100000010001010000100000001000100100110110",
--  (2058) iterative_modular_reduction_51
-- reg_a = o2_X; reg_b = prime2; reg_acc = reg_o >> 256; o2_X = reg_o; operation : s*b + a + acc
"000000100001100000010001010000100000001101001001010110",
--  (2059) iterative_modular_reduction_52
-- reg_a = o3_X; reg_b = prime3; reg_acc = reg_o >> 256; o3_X = reg_o; operation : s*b + a + acc
"000000100001100000010001010000100000010001101101110110",
--  (2060) iterative_modular_reduction_53
-- reg_a = o4_X; reg_b = prime4; reg_acc = reg_o >> 256; o4_X = reg_o; Enable sign a,b; operation : s*b + a + acc
"000000100001100000010001010000100001110110010010010110",
--  (2061) iterative_modular_reduction_54
-- NOP 4 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : b + a + acc;
"000000000000000100000000010000011110000100000000000010",
--  (2062) iterative_modular_reduction_55
-- -- In case of size 6
-- reg_a = a5_X; reg_b = 0; reg_acc = 0; Enable sign a,b; operation : b + a + acc;
"000000100001101000000000010000011001111010110110110010",
--  (2063) iterative_modular_reduction_56
-- reg_a = a0_X; reg_b = prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_positive; operation : -s*b + a + acc
"000000100001101000010011000111010000000100000000010010",
--  (2064) iterative_modular_reduction_57
-- reg_a = a1_X; reg_b = prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : -s*b + a + acc
"000000100001101000010011000000100000001000100100110010",
--  (2065) iterative_modular_reduction_58
-- reg_a = a2_X; reg_b = prime2; reg_acc = reg_o >> 256; o2_X = reg_o; operation : -s*b + a + acc
"000000100001101000010011000000100000001101001001010010",
--  (2066) iterative_modular_reduction_59
-- reg_a = a3_X; reg_b = prime3; reg_acc = reg_o >> 256; o3_X = reg_o; operation : -s*b + a + acc
"000000100001101000010011000000100000010001101101110010",
--  (2067) iterative_modular_reduction_60
-- reg_a = a4_X; reg_b = prime4; reg_acc = reg_o >> 256; o4_X = reg_o; operation : -s*b + a + acc
"000000100001101000010011000000100000010110010010010010",
--  (2068) iterative_modular_reduction_61
-- reg_a = a5_X; reg_b = prime5; reg_acc = reg_o >> 256; o5_X = reg_o; Enable sign a,b; operation : -s*b + a + acc
"000000100001101000010011000000100001111010110110110010",
--  (2069) iterative_modular_reduction_62
-- reg_a = o0_X; reg_b = prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc
"000000100001101000010001010011010000000100000000010110",
--  (2070) iterative_modular_reduction_63
-- reg_a = o1_X; reg_b = prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : s*b + a + acc
"000000100001101000010001010000100000001000100100110110",
--  (2071) iterative_modular_reduction_64
-- reg_a = o2_X; reg_b = prime2; reg_acc = reg_o >> 256; o2_X = reg_o; operation : s*b + a + acc
"000000100001101000010001010000100000001101001001010110",
--  (2072) iterative_modular_reduction_65
-- reg_a = o3_X; reg_b = prime3; reg_acc = reg_o >> 256; o3_X = reg_o; operation : s*b + a + acc
"000000100001101000010001010000100000010001101101110110",
--  (2073) iterative_modular_reduction_66
-- reg_a = o4_X; reg_b = prime4; reg_acc = reg_o >> 256; o4_X = reg_o; operation : s*b + a + acc
"000000100001101000010001010000100000010110010010010110",
--  (2074) iterative_modular_reduction_67
-- reg_a = o5_X; reg_b = prime5; reg_acc = reg_o >> 256; o5_X = reg_o; Enable sign a,b; operation : s*b + a + acc
"000000100001101000010001010000100001111010110110110110",
--  (2075) iterative_modular_reduction_68
-- reg_a = o0_X; reg_b = prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc
"000000100001101000010001010011010000000100000000010110",
--  (2076) iterative_modular_reduction_69
-- reg_a = o1_X; reg_b = prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : s*b + a + acc
"000000100001101000010001010000100000001000100100110110",
--  (2077) iterative_modular_reduction_70
-- reg_a = o2_X; reg_b = prime2; reg_acc = reg_o >> 256; o2_X = reg_o; operation : s*b + a + acc
"000000100001101000010001010000100000001101001001010110",
--  (2078) iterative_modular_reduction_71
-- reg_a = o3_X; reg_b = prime3; reg_acc = reg_o >> 256; o3_X = reg_o; operation : s*b + a + acc
"000000100001101000010001010000100000010001101101110110",
--  (2079) iterative_modular_reduction_72
-- reg_a = o4_X; reg_b = prime4; reg_acc = reg_o >> 256; o4_X = reg_o; operation : s*b + a + acc
"000000100001101000010001010000100000010110010010010110",
--  (2080) iterative_modular_reduction_73
-- reg_a = o5_X; reg_b = prime5; reg_acc = reg_o >> 256; o5_X = reg_o; Enable sign a,b; operation : s*b + a + acc
"000000100001101000010001010000100001111010110110110110",
--  (2081) iterative_modular_reduction_74
-- NOP 4 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : b + a + acc;
"000000000000000100000000010000011110000100000000000010",
--  (2082) iterative_modular_reduction_75
-- -- In case of size 7
-- reg_a = a6_X; reg_b = 0; reg_acc = 0; Enable sign a,b; operation : b + a + acc;
"000000100001110000000000010000011001111111011011010010",
--  (2083) iterative_modular_reduction_76
-- reg_a = a0_X; reg_b = prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_positive; operation : -s*b + a + acc
"000000100001110000010011000111010000000100000000010010",
--  (2084) iterative_modular_reduction_77
-- reg_a = a1_X; reg_b = prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : -s*b + a + acc
"000000100001110000010011000000100000001000100100110010",
--  (2085) iterative_modular_reduction_78
-- reg_a = a2_X; reg_b = prime2; reg_acc = reg_o >> 256; o2_X = reg_o; operation : -s*b + a + acc
"000000100001110000010011000000100000001101001001010010",
--  (2086) iterative_modular_reduction_79
-- reg_a = a3_X; reg_b = prime3; reg_acc = reg_o >> 256; o3_X = reg_o; operation : -s*b + a + acc
"000000100001110000010011000000100000010001101101110010",
--  (2087) iterative_modular_reduction_80
-- reg_a = a4_X; reg_b = prime4; reg_acc = reg_o >> 256; o4_X = reg_o; operation : -s*b + a + acc
"000000100001110000010011000000100000010110010010010010",
--  (2088) iterative_modular_reduction_81
-- reg_a = a5_X; reg_b = prime5; reg_acc = reg_o >> 256; o5_X = reg_o; operation : -s*b + a + acc
"000000100001110000010011000000100000011010110110110010",
--  (2089) iterative_modular_reduction_82
-- reg_a = a6_X; reg_b = prime6; reg_acc = reg_o >> 256; o6_X = reg_o; Enable sign a,b; operation : -s*b + a + acc
"000000100001110000010011000000100001111111011011010010",
--  (2090) iterative_modular_reduction_83
-- reg_a = o0_X; reg_b = prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc
"000000100001110000010001010011010000000100000000010110",
--  (2091) iterative_modular_reduction_84
-- reg_a = o1_X; reg_b = prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : s*b + a + acc
"000000100001110000010001010000100000001000100100110110",
--  (2092) iterative_modular_reduction_85
-- reg_a = o2_X; reg_b = prime2; reg_acc = reg_o >> 256; o2_X = reg_o; operation : s*b + a + acc
"000000100001110000010001010000100000001101001001010110",
--  (2093) iterative_modular_reduction_86
-- reg_a = o3_X; reg_b = prime3; reg_acc = reg_o >> 256; o3_X = reg_o; operation : s*b + a + acc
"000000100001110000010001010000100000010001101101110110",
--  (2094) iterative_modular_reduction_87
-- reg_a = o4_X; reg_b = prime4; reg_acc = reg_o >> 256; o4_X = reg_o; operation : s*b + a + acc
"000000100001110000010001010000100000010110010010010110",
--  (2095) iterative_modular_reduction_88
-- reg_a = o5_X; reg_b = prime5; reg_acc = reg_o >> 256; o5_X = reg_o; operation : s*b + a + acc
"000000100001110000010001010000100000011010110110110110",
--  (2096) iterative_modular_reduction_89
-- reg_a = o6_X; reg_b = prime6; reg_acc = reg_o >> 256; o6_X = reg_o; Enable sign a,b; operation : s*b + a + acc
"000000100001110000010001010000100001111111011011010110",
--  (2097) iterative_modular_reduction_90
-- reg_a = o0_X; reg_b = prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc
"000000100001110000010001010011010000000100000000010110",
--  (2098) iterative_modular_reduction_91
-- reg_a = o1_X; reg_b = prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : s*b + a + acc
"000000100001110000010001010000100000001000100100110110",
--  (2099) iterative_modular_reduction_92
-- reg_a = o2_X; reg_b = prime2; reg_acc = reg_o >> 256; o2_X = reg_o; operation : s*b + a + acc
"000000100001110000010001010000100000001101001001010110",
--  (2100) iterative_modular_reduction_93
-- reg_a = o3_X; reg_b = prime3; reg_acc = reg_o >> 256; o3_X = reg_o; operation : s*b + a + acc
"000000100001110000010001010000100000010001101101110110",
--  (2101) iterative_modular_reduction_94
-- reg_a = o4_X; reg_b = prime4; reg_acc = reg_o >> 256; o4_X = reg_o; operation : s*b + a + acc
"000000100001110000010001010000100000010110010010010110",
--  (2102) iterative_modular_reduction_95
-- reg_a = o5_X; reg_b = prime5; reg_acc = reg_o >> 256; o5_X = reg_o; operation : s*b + a + acc
"000000100001110000010001010000100000011010110110110110",
--  (2103) iterative_modular_reduction_96
-- reg_a = o6_X; reg_b = prime6; reg_acc = reg_o >> 256; o6_X = reg_o; Enable sign a,b; operation : s*b + a + acc
"000000100001110000010001010000100001111111011011010110",
--  (2104) iterative_modular_reduction_97
-- NOP 4 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : b + a + acc;
"000000000000000100000000010000011110000100000000000010",
--  (2105) iterative_modular_reduction_98
-- -- In case of size 8
-- reg_a = a7_X; reg_b = 0; reg_acc = 0; Enable sign a,b; operation : b + a + acc;
"000000100001111000000000010000011001100011111111110010",
--  (2106) iterative_modular_reduction_99
-- reg_a = a0_X; reg_b = prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_positive; operation : -s*b + a + acc
"000000100001111000010011000111010000000100000000010010",
--  (2107) iterative_modular_reduction_100
-- reg_a = a1_X; reg_b = prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : -s*b + a + acc
"000000100001111000010011000000100000001000100100110010",
--  (2108) iterative_modular_reduction_101
-- reg_a = a2_X; reg_b = prime2; reg_acc = reg_o >> 256; o2_X = reg_o; operation : -s*b + a + acc
"000000100001111000010011000000100000001101001001010010",
--  (2109) iterative_modular_reduction_102
-- reg_a = a3_X; reg_b = prime3; reg_acc = reg_o >> 256; o3_X = reg_o; operation : -s*b + a + acc
"000000100001111000010011000000100000010001101101110010",
--  (2110) iterative_modular_reduction_103
-- reg_a = a4_X; reg_b = prime4; reg_acc = reg_o >> 256; o4_X = reg_o; operation : -s*b + a + acc
"000000100001111000010011000000100000010110010010010010",
--  (2111) iterative_modular_reduction_104
-- reg_a = a5_X; reg_b = prime5; reg_acc = reg_o >> 256; o5_X = reg_o; operation : -s*b + a + acc
"000000100001111000010011000000100000011010110110110010",
--  (2112) iterative_modular_reduction_105
-- reg_a = a6_X; reg_b = prime6; reg_acc = reg_o >> 256; o6_X = reg_o; operation : -s*b + a + acc
"000000100001111000010011000000100000011111011011010010",
--  (2113) iterative_modular_reduction_106
-- reg_a = a7_X; reg_b = prime7; reg_acc = reg_o >> 256; o7_X = reg_o; Enable sign a,b; operation : -s*b + a + acc
"000000100001111000010011000000100001100011111111110010",
--  (2114) iterative_modular_reduction_107
-- reg_a = o0_X; reg_b = prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc
"000000100001111000010001010011010000000100000000010110",
--  (2115) iterative_modular_reduction_108
-- reg_a = o1_X; reg_b = prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : s*b + a + acc
"000000100001111000010001010000100000001000100100110110",
--  (2116) iterative_modular_reduction_109
-- reg_a = o2_X; reg_b = prime2; reg_acc = reg_o >> 256; o2_X = reg_o; operation : s*b + a + acc
"000000100001111000010001010000100000001101001001010110",
--  (2117) iterative_modular_reduction_110
-- reg_a = o3_X; reg_b = prime3; reg_acc = reg_o >> 256; o3_X = reg_o; operation : s*b + a + acc
"000000100001111000010001010000100000010001101101110110",
--  (2118) iterative_modular_reduction_111
-- reg_a = o4_X; reg_b = prime4; reg_acc = reg_o >> 256; o4_X = reg_o; operation : s*b + a + acc
"000000100001111000010001010000100000010110010010010110",
--  (2119) iterative_modular_reduction_112
-- reg_a = o5_X; reg_b = prime5; reg_acc = reg_o >> 256; o5_X = reg_o; operation : s*b + a + acc
"000000100001111000010001010000100000011010110110110110",
--  (2120) iterative_modular_reduction_113
-- reg_a = o6_X; reg_b = prime6; reg_acc = reg_o >> 256; o6_X = reg_o; operation : s*b + a + acc
"000000100001111000010001010000100000011111011011010110",
--  (2121) iterative_modular_reduction_114
-- reg_a = o7_X; reg_b = prime7; reg_acc = reg_o >> 256; o7_X = reg_o; Enable sign a,b; operation : s*b + a + acc
"000000100001111000010001010000100001100011111111110110",
--  (2122) iterative_modular_reduction_115
-- reg_a = o0_X; reg_b = prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc
"000000100001111000010001010011010000000100000000010110",
--  (2123) iterative_modular_reduction_116
-- reg_a = o1_X; reg_b = prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : s*b + a + acc
"000000100001111000010001010000100000001000100100110110",
--  (2124) iterative_modular_reduction_117
-- reg_a = o2_X; reg_b = prime2; reg_acc = reg_o >> 256; o2_X = reg_o; operation : s*b + a + acc
"000000100001111000010001010000100000001101001001010110",
--  (2125) iterative_modular_reduction_118
-- reg_a = o3_X; reg_b = prime3; reg_acc = reg_o >> 256; o3_X = reg_o; operation : s*b + a + acc
"000000100001111000010001010000100000010001101101110110",
--  (2126) iterative_modular_reduction_119
-- reg_a = o4_X; reg_b = prime4; reg_acc = reg_o >> 256; o4_X = reg_o; operation : s*b + a + acc
"000000100001111000010001010000100000010110010010010110",
--  (2127) iterative_modular_reduction_120
-- reg_a = o5_X; reg_b = prime5; reg_acc = reg_o >> 256; o5_X = reg_o; operation : s*b + a + acc
"000000100001111000010001010000100000011010110110110110",
--  (2128) iterative_modular_reduction_121
-- reg_a = o6_X; reg_b = prime6; reg_acc = reg_o >> 256; o6_X = reg_o; operation : s*b + a + acc
"000000100001111000010001010000100000011111011011010110",
--  (2129) iterative_modular_reduction_122
-- reg_a = o7_X; reg_b = prime7; reg_acc = reg_o >> 256; o7_X = reg_o; Enable sign a,b; operation : s*b + a + acc
"000000100001111000010001010000100001100011111111110110",
--  (2130) iterative_modular_reduction_123
-- NOP 4 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : b + a + acc;
"000000000000000100000000010000011110000100000000000010",
--  (2131) addition_subtraction_with_reduction_0
-- Operands size 1
-- reg_a = a0_X; reg_b = b0_X; reg_acc = 0; o0_X = reg_o; Enable sign a,b; operation : b +/- a + acc;
"000000100001000000010000011000010001100100000000000010",
--  (2132) addition_subtraction_with_reduction_1
-- reg_a = 0; reg_b = 2prime0; reg_acc = reg_o; reg_s = reg_o_positive; o0_X = reg_o; Enable sign a,b; operation : -s*b + a + acc;
"000000100001000000010011000111000111100100000000001010",
--  (2133) addition_subtraction_with_reduction_2
-- reg_a = 0; reg_b = 2prime0; reg_acc = reg_o; reg_s = reg_o_negative; o0_X = reg_o; Enable sign a,b; operation : s*b + a + acc;
"000000100001000000010001010011000111100100000000001010",
--  (2134) addition_subtraction_with_reduction_3
-- reg_a = 0; reg_b = 2prime0; reg_acc = reg_o; reg_s = reg_o_negative; o0_X = reg_o; Enable sign a,b; operation : s*b + a + acc;
"000000100001000000010001010011000111100100000000001010",
--  (2135) addition_subtraction_with_reduction_4
-- NOP 4 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : b + a + acc;
"000000000000000100000000010000011110000100000000000010",
--  (2136) addition_subtraction_with_reduction_5
-- -- In case of sizes 2, 3, 4, 5, 6, 7, 8
-- reg_a = a0_X; reg_b = b0_X; reg_acc = 0; o0_X = reg_o; operation : b +/- a + acc;
"000100100001001000010000001000010000000100000000000010",
--  (2137) addition_subtraction_with_reduction_6
-- -- In case of size 2
-- reg_a = a1_X; reg_b = b1_X; reg_acc = reg_o >> 256; o1_X = reg_o; Enable sign a, b; operation : b +/- a + acc;
"000000100001001000010000001000100001101000100100100010",
--  (2138) addition_subtraction_with_reduction_7
-- reg_a = o0_X; reg_b = 2prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_positive; operation : -s*b + a + acc;
"000000100001001000010011000111010000000100000000001110",
--  (2139) addition_subtraction_with_reduction_8
-- reg_a = o1_X; reg_b = 2prime1; reg_acc = reg_o >> 256; o1_X = reg_o; Enable sign a,b; operation : -s*b + a + acc;
"000000100001001000010011000000100001101000100100101110",
--  (2140) addition_subtraction_with_reduction_9
-- reg_a = o0_X; reg_b = 2prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc;
"000000100001001000010001010011010000000100000000001110",
--  (2141) addition_subtraction_with_reduction_10
-- reg_a = o1_X; reg_b = 2prime1; reg_acc = reg_o >> 256; o1_X = reg_o; Enable sign a,b; operation : s*b + a + acc;
"000000100001001000010001010000100001101000100100101110",
--  (2142) addition_subtraction_with_reduction_11
-- reg_a = o0_X; reg_b = 2prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc;
"000000100001001000010001010011010000000100000000001110",
--  (2143) addition_subtraction_with_reduction_12
-- reg_a = o1_X; reg_b = 2prime1; reg_acc = reg_o >> 256; o1_X = reg_o; Enable sign a,b; operation : s*b + a + acc;
"000000100001001000010001010000100001101000100100101110",
--  (2144) addition_subtraction_with_reduction_13
-- NOP 4 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : b + a + acc;
"000000000000000100000000010000011110000100000000000010",
--  (2145) addition_subtraction_with_reduction_14
-- -- In case of sizes 3, 4, 5, 6, 7, 8
-- reg_a = a1_X; reg_b = b1_X; reg_acc = reg_o >> 256; o1_X = reg_o; operation : b +/- a + acc;
"000110000001010000010000001000100000001000100100100010",
--  (2146) addition_subtraction_with_reduction_15
-- -- In case of size 3
-- reg_a = a2_X; reg_b = b2_X; reg_acc = reg_o >> 256; o2_X = reg_o; Enable sign a, b; operation : b +/- a + acc;
"000000100001010000010000001000100001100101001001000010",
--  (2147) addition_subtraction_with_reduction_16
-- reg_a = o0_X; reg_b = 2prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_positive; operation : -s*b + a + acc;
"000000100001010000010011000111010000000100000000001110",
--  (2148) addition_subtraction_with_reduction_17
-- reg_a = o1_X; reg_b = 2prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : -s*b + a + acc;
"000000100001010000010011000000100000001000100100101110",
--  (2149) addition_subtraction_with_reduction_18
-- reg_a = o2_X; reg_b = 2prime2; reg_acc = reg_o >> 256; o2_X = reg_o; Enable sign a,b; operation : -s*b + a + acc;
"000000100001010000010011000000100001101101001001001110",
--  (2150) addition_subtraction_with_reduction_19
-- reg_a = o0_X; reg_b = 2prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc;
"000000100001010000010001010011010000000100000000001110",
--  (2151) addition_subtraction_with_reduction_20
-- reg_a = o1_X; reg_b = 2prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : s*b + a + acc;
"000000100001010000010001010000100000001000100100101110",
--  (2152) addition_subtraction_with_reduction_21
-- reg_a = o2_X; reg_b = 2prime2; reg_acc = reg_o >> 256; o2_X = reg_o; Enable sign a,b; operation : s*b + a + acc;
"000000100001010000010001010000100001101101001001001110",
--  (2153) addition_subtraction_with_reduction_22
-- reg_a = o0_X; reg_b = 2prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc;
"000000100001010000010001010011010000000100000000001110",
--  (2154) addition_subtraction_with_reduction_23
-- reg_a = o1_X; reg_b = 2prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : s*b + a + acc;
"000000100001010000010001010000100000001000100100101110",
--  (2155) addition_subtraction_with_reduction_24
-- reg_a = o2_X; reg_b = 2prime2; reg_acc = reg_o >> 256; o2_X = reg_o; Enable sign a,b; operation : s*b + a + acc;
"000000100001010000010001010000100001101101001001001110",
--  (2156) addition_subtraction_with_reduction_25
-- NOP 4 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : b + a + acc;
"000000000000000100000000010000011110000100000000000010",
--  (2157) addition_subtraction_with_reduction_26
-- -- In case of size 4, 5, 6, 7, 8
-- reg_a = a2_X; reg_b = b2_X; reg_acc = reg_o >> 256; o2_X = reg_o; operation : b +/- a + acc;
"000111100001011000010000001000100000000101001001000010",
--  (2158) addition_subtraction_with_reduction_27
-- -- In case of size 4
-- reg_a = a3_X; reg_b = b3_X; reg_acc = reg_o >> 256; o3_X = reg_o; Enable sign a, b; operation : b +/- a + acc;
"000000100001011000010000001000100001110001101101100010",
--  (2159) addition_subtraction_with_reduction_28
-- reg_a = o0_X; reg_b = 2prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_positive; operation : -s*b + a + acc;
"000000100001011000010011000111010000000100000000001110",
--  (2160) addition_subtraction_with_reduction_29
-- reg_a = o1_X; reg_b = 2prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : -s*b + a + acc;
"000000100001011000010011000000100000001000100100101110",
--  (2161) addition_subtraction_with_reduction_30
-- reg_a = o2_X; reg_b = 2prime2; reg_acc = reg_o >> 256; o2_X = reg_o; operation : -s*b + a + acc;
"000000100001011000010011000000100000001101001001001110",
--  (2162) addition_subtraction_with_reduction_31
-- reg_a = o3_X; reg_b = 2prime3; reg_acc = reg_o >> 256; o3_X = reg_o; Enable sign a,b; operation : -s*b + a + acc;
"000000100001011000010011000000100001100001101101101110",
--  (2163) addition_subtraction_with_reduction_32
-- reg_a = o0_X; reg_b = 2prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc;
"000000100001011000010001010011010000000100000000001110",
--  (2164) addition_subtraction_with_reduction_33
-- reg_a = o1_X; reg_b = 2prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : s*b + a + acc;
"000000100001011000010001010000100000001000100100101110",
--  (2165) addition_subtraction_with_reduction_34
-- reg_a = o2_X; reg_b = 2prime2; reg_acc = reg_o >> 256; o2_X = reg_o; operation : s*b + a + acc;
"000000100001011000010001010000100000001101001001001110",
--  (2166) addition_subtraction_with_reduction_35
-- reg_a = o3_X; reg_b = 2prime3; reg_acc = reg_o >> 256; o3_X = reg_o; Enable sign a,b; operation : s*b + a + acc;
"000000100001011000010001010000100001100001101101101110",
--  (2167) addition_subtraction_with_reduction_36
-- reg_a = o0_X; reg_b = 2prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc;
"000000100001011000010001010011010000000100000000001110",
--  (2168) addition_subtraction_with_reduction_37
-- reg_a = o1_X; reg_b = 2prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : s*b + a + acc;
"000000100001011000010001010000100000001000100100101110",
--  (2169) addition_subtraction_with_reduction_38
-- reg_a = o2_X; reg_b = 2prime2; reg_acc = reg_o >> 256; o2_X = reg_o; operation : s*b + a + acc;
"000000100001011000010001010000100000001101001001001110",
--  (2170) addition_subtraction_with_reduction_39
-- reg_a = o3_X; reg_b = 2prime3; reg_acc = reg_o >> 256; o3_X = reg_o; Enable sign a,b; operation : s*b + a + acc;
"000000100001011000010001010000100001110001101101101110",
--  (2171) addition_subtraction_with_reduction_40
-- NOP 4 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : b + a + acc;
"000000000000000100000000010000011110000100000000000010",
--  (2172) addition_subtraction_with_reduction_41
-- -- In case of size 5, 6, 7, 8
-- reg_a = a3_X; reg_b = b3_X; reg_acc = reg_o >> 256; o3_X = reg_o; operation : b +/- a + acc;
"001001000001100000010000001000100000010001101101100010",
--  (2173) addition_subtraction_with_reduction_42
-- -- In case of size 5
-- reg_a = a4_X; reg_b = b4_X; reg_acc = reg_o >> 256; o4_X = reg_o; Enable sign a, b; operation : b +/- a + acc;
"000000100001100000010000001000100001110110010010000010",
--  (2174) addition_subtraction_with_reduction_43
-- reg_a = o0_X; reg_b = 2prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_positive; operation : -s*b + a + acc;
"000000100001100000010011000111010000000100000000001110",
--  (2175) addition_subtraction_with_reduction_44
-- reg_a = o1_X; reg_b = 2prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : -s*b + a + acc;
"000000100001100000010011000000100000001000100100101110",
--  (2176) addition_subtraction_with_reduction_45
-- reg_a = o2_X; reg_b = 2prime2; reg_acc = reg_o >> 256; o2_X = reg_o; operation : -s*b + a + acc;
"000000100001100000010011000000100000001101001001001110",
--  (2177) addition_subtraction_with_reduction_46
-- reg_a = o3_X; reg_b = 2prime3; reg_acc = reg_o >> 256; o3_X = reg_o; operation : -s*b + a + acc;
"000000100001100000010011000000100000010001101101101110",
--  (2178) addition_subtraction_with_reduction_47
-- reg_a = o4_X; reg_b = 2prime4; reg_acc = reg_o >> 256; o4_X = reg_o; Enable sign a,b; operation : -s*b + a + acc;
"000000100001100000010011000000100001110110010010001110",
--  (2179) addition_subtraction_with_reduction_48
-- reg_a = o0_X; reg_b = 2prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc;
"000000100001100000010001010011010000000100000000001110",
--  (2180) addition_subtraction_with_reduction_49
-- reg_a = o1_X; reg_b = 2prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : s*b + a + acc;
"000000100001100000010001010000100000001000100100101110",
--  (2181) addition_subtraction_with_reduction_50
-- reg_a = o2_X; reg_b = 2prime2; reg_acc = reg_o >> 256; o2_X = reg_o; operation : s*b + a + acc;
"000000100001100000010001010000100000001101001001001110",
--  (2182) addition_subtraction_with_reduction_51
-- reg_a = o3_X; reg_b = 2prime3; reg_acc = reg_o >> 256; o3_X = reg_o; operation : s*b + a + acc;
"000000100001100000010001010000100000010001101101101110",
--  (2183) addition_subtraction_with_reduction_52
-- reg_a = o4_X; reg_b = 2prime4; reg_acc = reg_o >> 256; o4_X = reg_o; Enable sign a,b; operation : s*b + a + acc;
"000000100001100000010001010000100001110110010010001110",
--  (2184) addition_subtraction_with_reduction_53
-- reg_a = o0_X; reg_b = 2prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc;
"000000100001100000010001010011010000000100000000001110",
--  (2185) addition_subtraction_with_reduction_54
-- reg_a = o1_X; reg_b = 2prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : s*b + a + acc;
"000000100001100000010001010000100000001000100100101110",
--  (2186) addition_subtraction_with_reduction_55
-- reg_a = o2_X; reg_b = 2prime2; reg_acc = reg_o >> 256; o2_X = reg_o; operation : s*b + a + acc;
"000000100001100000010001010000100000001101001001001110",
--  (2187) addition_subtraction_with_reduction_56
-- reg_a = o3_X; reg_b = 2prime3; reg_acc = reg_o >> 256; o3_X = reg_o; operation : s*b + a + acc;
"000000100001100000010001010000100000010001101101101110",
--  (2188) addition_subtraction_with_reduction_57
-- reg_a = o4_X; reg_b = 2prime4; reg_acc = reg_o >> 256; o4_X = reg_o; Enable sign a,b; operation : s*b + a + acc;
"000000100001100000010001010000100001110110010010001110",
--  (2189) addition_subtraction_with_reduction_58
-- NOP 4 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : b + a + acc;
"000000000000000100000000010000011110000100000000000010",
--  (2190) addition_subtraction_with_reduction_59
-- -- In case of size 6, 7, 8
-- reg_a = a4_X; reg_b = b4_X; reg_acc = reg_o >> 256; o4_X = reg_o; operation : b +/- a + acc;
"001010100001101000010000001000100000010110010010000010",
--  (2191) addition_subtraction_with_reduction_60
-- -- In case of size 6
-- reg_a = a5_X; reg_b = b5_X; reg_acc = reg_o >> 256; o5_X = reg_o; Enable sign a, b; operation : b +/- a + acc;
"000000100001101000010000001000100001111010110110100010",
--  (2192) addition_subtraction_with_reduction_61
-- reg_a = o0_X; reg_b = 2prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_positive; operation : -s*b + a + acc;
"000000100001101000010011000111010000000100000000001110",
--  (2193) addition_subtraction_with_reduction_62
-- reg_a = o1_X; reg_b = 2prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : -s*b + a + acc;
"000000100001101000010011000000100000001000100100101110",
--  (2194) addition_subtraction_with_reduction_63
-- reg_a = o2_X; reg_b = 2prime2; reg_acc = reg_o >> 256; o2_X = reg_o; operation : -s*b + a + acc;
"000000100001101000010011000000100000001101001001001110",
--  (2195) addition_subtraction_with_reduction_64
-- reg_a = o3_X; reg_b = 2prime3; reg_acc = reg_o >> 256; o3_X = reg_o; operation : -s*b + a + acc;
"000000100001101000010011000000100000010001101101101110",
--  (2196) addition_subtraction_with_reduction_65
-- reg_a = o4_X; reg_b = 2prime4; reg_acc = reg_o >> 256; o4_X = reg_o; operation : -s*b + a + acc;
"000000100001101000010011000000100000010110010010001110",
--  (2197) addition_subtraction_with_reduction_66
-- reg_a = o5_X; reg_b = 2prime5; reg_acc = reg_o >> 256; o5_X = reg_o; Enable sign a,b; operation : -s*b + a + acc;
"000000100001101000010011000000100001111010110110101110",
--  (2198) addition_subtraction_with_reduction_67
-- reg_a = o0_X; reg_b = 2prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc;
"000000100001101000010001010011010000000100000000001110",
--  (2199) addition_subtraction_with_reduction_68
-- reg_a = o1_X; reg_b = 2prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : s*b + a + acc;
"000000100001101000010001010000100000001000100100101110",
--  (2200) addition_subtraction_with_reduction_69
-- reg_a = o2_X; reg_b = 2prime2; reg_acc = reg_o >> 256; o2_X = reg_o; operation : s*b + a + acc;
"000000100001101000010001010000100000001101001001001110",
--  (2201) addition_subtraction_with_reduction_70
-- reg_a = o3_X; reg_b = 2prime3; reg_acc = reg_o >> 256; o3_X = reg_o; operation : s*b + a + acc;
"000000100001101000010001010000100000010001101101101110",
--  (2202) addition_subtraction_with_reduction_71
-- reg_a = o4_X; reg_b = 2prime4; reg_acc = reg_o >> 256; o4_X = reg_o; operation : s*b + a + acc;
"000000100001101000010001010000100000010110010010001110",
--  (2203) addition_subtraction_with_reduction_72
-- reg_a = o5_X; reg_b = 2prime5; reg_acc = reg_o >> 256; o5_X = reg_o; Enable sign a,b; operation : s*b + a + acc;
"000000100001101000010001010000100001111010110110101110",
--  (2204) addition_subtraction_with_reduction_73
-- reg_a = o0_X; reg_b = 2prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc;
"000000100001101000010001010011010000000100000000001110",
--  (2205) addition_subtraction_with_reduction_74
-- reg_a = o1_X; reg_b = 2prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : s*b + a + acc;
"000000100001101000010001010000100000001000100100101110",
--  (2206) addition_subtraction_with_reduction_75
-- reg_a = o2_X; reg_b = 2prime2; reg_acc = reg_o >> 256; o2_X = reg_o; operation : s*b + a + acc;
"000000100001101000010001010000100000001101001001001110",
--  (2207) addition_subtraction_with_reduction_76
-- reg_a = o3_X; reg_b = 2prime3; reg_acc = reg_o >> 256; o3_X = reg_o; operation : s*b + a + acc;
"000000100001101000010001010000100000010001101101101110",
--  (2208) addition_subtraction_with_reduction_77
-- reg_a = o4_X; reg_b = 2prime4; reg_acc = reg_o >> 256; o4_X = reg_o; operation : s*b + a + acc;
"000000100001101000010001010000100000010110010010001110",
--  (2209) addition_subtraction_with_reduction_78
-- reg_a = o5_X; reg_b = 2prime5; reg_acc = reg_o >> 256; o5_X = reg_o; Enable sign a,b; operation : s*b + a + acc;
"000000100001101000010001010000100001111010110110101110",
--  (2210) addition_subtraction_with_reduction_79
-- NOP 4 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : b + a + acc;
"000000000000000100000000010000011110000100000000000010",
--  (2211) addition_subtraction_with_reduction_80
-- -- In case of size 7, 8
-- reg_a = a5_X; reg_b = b5_X; reg_acc = reg_o >> 256; o5_X = reg_o; operation : b +/- a + acc;
"001100000001110000010000001000100000011010110110100010",
--  (2212) addition_subtraction_with_reduction_81
-- -- In case of size 7
-- reg_a = a6_X; reg_b = b6_X; reg_acc = reg_o >> 256; o6_X = reg_o; Enable sign a, b; operation : b +/- a + acc;
"000000100001110000010000001000100001111111011011000010",
--  (2213) addition_subtraction_with_reduction_82
-- reg_a = o0_X; reg_b = 2prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_positive; operation : -s*b + a + acc;
"000000100001110000010011000111010000000100000000001110",
--  (2214) addition_subtraction_with_reduction_83
-- reg_a = o1_X; reg_b = 2prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : -s*b + a + acc;
"000000100001110000010011000000100000001000100100101110",
--  (2215) addition_subtraction_with_reduction_84
-- reg_a = o2_X; reg_b = 2prime2; reg_acc = reg_o >> 256; o2_X = reg_o; operation : -s*b + a + acc;
"000000100001110000010011000000100000001101001001001110",
--  (2216) addition_subtraction_with_reduction_85
-- reg_a = o3_X; reg_b = 2prime3; reg_acc = reg_o >> 256; o3_X = reg_o; operation : -s*b + a + acc;
"000000100001110000010011000000100000010001101101101110",
--  (2217) addition_subtraction_with_reduction_86
-- reg_a = o4_X; reg_b = 2prime4; reg_acc = reg_o >> 256; o4_X = reg_o; operation : -s*b + a + acc;
"000000100001110000010011000000100000010110010010001110",
--  (2218) addition_subtraction_with_reduction_87
-- reg_a = o5_X; reg_b = 2prime5; reg_acc = reg_o >> 256; o5_X = reg_o; operation : -s*b + a + acc;
"000000100001110000010011000000100000011010110110101110",
--  (2219) addition_subtraction_with_reduction_88
-- reg_a = o6_X; reg_b = 2prime6; reg_acc = reg_o >> 256; o6_X = reg_o; Enable sign a,b; operation : -s*b + a + acc;
"000000100001110000010011000000100001111111011011001110",
--  (2220) addition_subtraction_with_reduction_89
-- reg_a = o0_X; reg_b = 2prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc;
"000000100001110000010001010011010000000100000000001110",
--  (2221) addition_subtraction_with_reduction_90
-- reg_a = o1_X; reg_b = 2prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : s*b + a + acc;
"000000100001110000010001010000100000001000100100101110",
--  (2222) addition_subtraction_with_reduction_91
-- reg_a = o2_X; reg_b = 2prime2; reg_acc = reg_o >> 256; o2_X = reg_o; operation : s*b + a + acc;
"000000100001110000010001010000100000001101001001001110",
--  (2223) addition_subtraction_with_reduction_92
-- reg_a = o3_X; reg_b = 2prime3; reg_acc = reg_o >> 256; o3_X = reg_o; operation : s*b + a + acc;
"000000100001110000010001010000100000010001101101101110",
--  (2224) addition_subtraction_with_reduction_93
-- reg_a = o4_X; reg_b = 2prime4; reg_acc = reg_o >> 256; o4_X = reg_o; operation : s*b + a + acc;
"000000100001110000010001010000100000010110010010001110",
--  (2225) addition_subtraction_with_reduction_94
-- reg_a = o5_X; reg_b = 2prime5; reg_acc = reg_o >> 256; o5_X = reg_o; operation : s*b + a + acc;
"000000100001110000010001010000100000011010110110101110",
--  (2226) addition_subtraction_with_reduction_95
-- reg_a = o6_X; reg_b = 2prime6; reg_acc = reg_o >> 256; o6_X = reg_o; Enable sign a,b; operation : s*b + a + acc;
"000000100001110000010001010000100001111111011011001110",
--  (2227) addition_subtraction_with_reduction_96
-- reg_a = o0_X; reg_b = 2prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc;
"000000100001110000010001010011010000000100000000001110",
--  (2228) addition_subtraction_with_reduction_97
-- reg_a = o1_X; reg_b = 2prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : s*b + a + acc;
"000000100001110000010001010000100000001000100100101110",
--  (2229) addition_subtraction_with_reduction_98
-- reg_a = o2_X; reg_b = 2prime2; reg_acc = reg_o >> 256; o2_X = reg_o; operation : s*b + a + acc;
"000000100001110000010001010000100000001101001001001110",
--  (2230) addition_subtraction_with_reduction_99
-- reg_a = o3_X; reg_b = 2prime3; reg_acc = reg_o >> 256; o3_X = reg_o; operation : s*b + a + acc;
"000000100001110000010001010000100000010001101101101110",
--  (2231) addition_subtraction_with_reduction_100
-- reg_a = o4_X; reg_b = 2prime4; reg_acc = reg_o >> 256; o4_X = reg_o; operation : s*b + a + acc;
"000000100001110000010001010000100000010110010010001110",
--  (2232) addition_subtraction_with_reduction_101
-- reg_a = o5_X; reg_b = 2prime5; reg_acc = reg_o >> 256; o5_X = reg_o; operation : s*b + a + acc;
"000000100001110000010001010000100000011010110110101110",
--  (2233) addition_subtraction_with_reduction_102
-- reg_a = o6_X; reg_b = 2prime6; reg_acc = reg_o >> 256; o6_X = reg_o; Enable sign a,b; operation : s*b + a + acc;
"000000100001110000010001010000100001111111011011001110",
--  (2234) addition_subtraction_with_reduction_103
-- NOP 4 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : b + a + acc;
"000000000000000100000000010000011110000100000000000010",
--  (2235) addition_subtraction_with_reduction_104
-- -- In case of size 8
-- reg_a = a6_X; reg_b = b6_X; reg_acc = reg_o >> 256; o6_X = reg_o; operation : b +/- a + acc;
"000000100001111000010000001000100000011111011011000010",
--  (2236) addition_subtraction_with_reduction_105
-- reg_a = a7_X; reg_b = b7_X; reg_acc = reg_o >> 256; o7_X = reg_o; Enable sign a,b; operation : b +/- a + acc;
"000000100001111000010000001000100001100011111111100010",
--  (2237) addition_subtraction_with_reduction_106
-- reg_a = o0_X; reg_b = 2prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_positive; operation : -s*b + a + acc;
"000000100001111000010011000111010000000100000000001110",
--  (2238) addition_subtraction_with_reduction_107
-- reg_a = o1_X; reg_b = 2prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : -s*b + a + acc;
"000000100001111000010011000000100000001000100100101110",
--  (2239) addition_subtraction_with_reduction_108
-- reg_a = o2_X; reg_b = 2prime2; reg_acc = reg_o >> 256; o2_X = reg_o; operation : -s*b + a + acc;
"000000100001111000010011000000100000001101001001001110",
--  (2240) addition_subtraction_with_reduction_109
-- reg_a = o3_X; reg_b = 2prime3; reg_acc = reg_o >> 256; o3_X = reg_o; operation : -s*b + a + acc;
"000000100001111000010011000000100000010001101101101110",
--  (2241) addition_subtraction_with_reduction_110
-- reg_a = o4_X; reg_b = 2prime4; reg_acc = reg_o >> 256; o4_X = reg_o; operation : -s*b + a + acc;
"000000100001111000010011000000100000010110010010001110",
--  (2242) addition_subtraction_with_reduction_111
-- reg_a = o5_X; reg_b = 2prime5; reg_acc = reg_o >> 256; o5_X = reg_o; operation : -s*b + a + acc;
"000000100001111000010011000000100000011010110110101110",
--  (2243) addition_subtraction_with_reduction_112
-- reg_a = o6_X; reg_b = 2prime6; reg_acc = reg_o >> 256; o6_X = reg_o; operation : -s*b + a + acc;
"000000100001111000010011000000100000011111011011001110",
--  (2244) addition_subtraction_with_reduction_113
-- reg_a = o7_X; reg_b = 2prime7; reg_acc = reg_o >> 256; o7_X = reg_o; Enable sign a,b; operation : -s*b + a + acc;
"000000100001111000010011000000100001100011111111101110",
--  (2245) addition_subtraction_with_reduction_114
-- reg_a = o0_X; reg_b = 2prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc;
"000000100001111000010001010011010000000100000000001110",
--  (2246) addition_subtraction_with_reduction_115
-- reg_a = o1_X; reg_b = 2prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : s*b + a + acc;
"000000100001111000010001010000100000001000100100101110",
--  (2247) addition_subtraction_with_reduction_116
-- reg_a = o2_X; reg_b = 2prime2; reg_acc = reg_o >> 256; o2_X = reg_o; operation : s*b + a + acc;
"000000100001111000010001010000100000001101001001001110",
--  (2248) addition_subtraction_with_reduction_117
-- reg_a = o3_X; reg_b = 2prime3; reg_acc = reg_o >> 256; o3_X = reg_o; operation : s*b + a + acc;
"000000100001111000010001010000100000010001101101101110",
--  (2249) addition_subtraction_with_reduction_118
-- reg_a = o4_X; reg_b = 2prime4; reg_acc = reg_o >> 256; o4_X = reg_o; operation : s*b + a + acc;
"000000100001111000010001010000100000010110010010001101",
--  (2250) addition_subtraction_with_reduction_119
-- reg_a = o5_X; reg_b = 2prime5; reg_acc = reg_o >> 256; o5_X = reg_o; operation : s*b + a + acc;
"000000100001111000010001010000100000011010110110101110",
--  (2251) addition_subtraction_with_reduction_120
-- reg_a = o6_X; reg_b = 2prime6; reg_acc = reg_o >> 256; o6_X = reg_o; operation : s*b + a + acc;
"000000100001111000010001010000100000011111011011001110",
--  (2252) addition_subtraction_with_reduction_121
-- reg_a = o7_X; reg_b = 2prime7; reg_acc = reg_o >> 256; o7_X = reg_o; Enable sign a,b; operation : s*b + a + acc;
"000000100001111000010001010000100001100011111111101110",
--  (2253) addition_subtraction_with_reduction_122
-- reg_a = o0_X; reg_b = 2prime0; reg_acc = 0; o0_X = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc;
"000000100001111000010001010011010000000100000000001110",
--  (2254) addition_subtraction_with_reduction_123
-- reg_a = o1_X; reg_b = 2prime1; reg_acc = reg_o >> 256; o1_X = reg_o; operation : s*b + a + acc;
"000000100001111000010001010000100000001000100100101110",
--  (2255) addition_subtraction_with_reduction_124
-- reg_a = o2_X; reg_b = 2prime2; reg_acc = reg_o >> 256; o2_X = reg_o; operation : s*b + a + acc;
"000000100001111000010001010000100000001101001001001110",
--  (2256) addition_subtraction_with_reduction_125
-- reg_a = o3_X; reg_b = 2prime3; reg_acc = reg_o >> 256; o3_X = reg_o; operation : s*b + a + acc;
"000000100001111000010001010000100000010001101101101110",
--  (2257) addition_subtraction_with_reduction_126
-- reg_a = o4_X; reg_b = 2prime4; reg_acc = reg_o >> 256; o4_X = reg_o; operation : s*b + a + acc;
"000000100001111000010001010000100000010110010010001110",
--  (2258) addition_subtraction_with_reduction_127
-- reg_a = o5_X; reg_b = 2prime5; reg_acc = reg_o >> 256; o5_X = reg_o; operation : s*b + a + acc;
"000000100001111000010001010000100000011010110110101110",
--  (2259) addition_subtraction_with_reduction_128
-- reg_a = o6_X; reg_b = 2prime6; reg_acc = reg_o >> 256; o6_X = reg_o; operation : s*b + a + acc;
"000000100001111000010001010000100000011111011011001110",
--  (2260) addition_subtraction_with_reduction_129
-- reg_a = o7_X; reg_b = 2prime7; reg_acc = reg_o >> 256; o7_X = reg_o; Enable sign a,b; operation : s*b + a + acc;
"000000100001111000010001010000100001100011111111101110",
--  (2261) addition_subtraction_with_reduction_130
-- NOP 4 stages                  
-- reg_a = 0; reg_b = 0; reg_acc = 0; operation : b + a + acc;
"000000000000000100000000010000011110000100000000000010"
);





constant rom_state_machine_fill_nop : romtype(2262 to 4095) := (others => "000000000000000100000000100000011110000100000000000011");
constant rom_state_machine : romtype(0 to 4095) := rom_state_machine_program & rom_state_machine_fill_nop;

signal rom_state_machine_address : std_logic_vector(11 downto 0);
signal rom_state_machine_next_address : std_logic_vector(11 downto 0);
signal rom_state_machine_output : std_logic_vector(53 downto 0);

signal rom_sm_rotation_size : std_logic_vector(1 downto 0);
signal rom_sel_address_a : std_logic;
signal rom_sel_address_b_prime : std_logic_vector(1 downto 0);
signal rom_sm_specific_mac_address_a : std_logic_vector(2 downto 0);
signal rom_sm_specific_mac_address_b : std_logic_vector(2 downto 0);
signal rom_sm_specific_mac_address_o : std_logic_vector(2 downto 0);
signal rom_sm_specific_mac_next_address_o : std_logic_vector(2 downto 0);
signal rom_mac_enable_signed_a : std_logic;
signal rom_mac_enable_signed_b : std_logic;
signal rom_mac_sel_load_reg_a : std_logic_vector(1 downto 0);
signal rom_mac_clear_reg_b : std_logic;
signal rom_mac_clear_reg_acc : std_logic;
signal rom_mac_sel_shift_reg_o : std_logic;
signal rom_mac_enable_update_reg_s : std_logic;
signal rom_mac_sel_reg_s_reg_o_sign : std_logic;
signal rom_mac_reg_s_reg_o_positive : std_logic;
signal rom_sm_sign_a_mode : std_logic;
signal rom_sm_mac_operation_mode : std_logic_vector(1 downto 0);
signal rom_mac_enable_reg_s_mask : std_logic;
signal rom_mac_subtraction_reg_a_b : std_logic;
signal rom_mac_sel_multiply_two_a_b : std_logic;
signal rom_mac_sel_reg_y_output : std_logic;
signal rom_sm_mac_write_enable_output : std_logic;
signal rom_mac_memory_double_mode : std_logic;
signal rom_mac_memory_only_write_mode : std_logic;
signal rom_base_address_generator_o_increment_previous_address : std_logic;

signal rom_last_state : std_logic;
signal rom_current_operand_size : std_logic_vector(2 downto 0);
signal rom_next_operation_same_operand_size : std_logic_vector(4 downto 0);
signal rom_next_operation_different_operand_size : std_logic_vector(6 downto 0);

signal adder_a : unsigned(11 downto 0);
signal adder_b : unsigned(6 downto 0);
signal adder_o : unsigned(11 downto 0);

signal ultimate_instruction : std_logic;

signal internal_sel_output_rom : std_logic;
signal internal_update_rom_address : std_logic;
signal internal_sel_load_new_rom_address : std_logic;
signal internal_sm_rotation_size : std_logic_vector(1 downto 0);
signal internal_sm_circular_shift_enable : std_logic;
signal internal_sel_address_a : std_logic;
signal internal_sel_address_b_prime : std_logic_vector(1 downto 0);
signal internal_sm_specific_mac_address_a : std_logic_vector(2 downto 0);
signal internal_sm_specific_mac_address_b : std_logic_vector(2 downto 0);
signal internal_sm_specific_mac_address_o : std_logic_vector(2 downto 0);
signal internal_sm_specific_mac_next_address_o : std_logic_vector(2 downto 0);
signal internal_mac_enable_signed_a : std_logic;
signal internal_mac_enable_signed_b : std_logic;
signal internal_mac_sel_load_reg_a : std_logic_vector(1 downto 0);
signal internal_mac_clear_reg_b : std_logic;
signal internal_mac_clear_reg_acc : std_logic;
signal internal_mac_sel_shift_reg_o : std_logic;
signal internal_mac_enable_update_reg_s : std_logic;
signal internal_mac_sel_reg_s_reg_o_sign : std_logic;
signal internal_mac_reg_s_reg_o_positive : std_logic;
signal internal_sm_sign_a_mode : std_logic;
signal internal_sm_mac_operation_mode : std_logic_vector(1 downto 0);
signal internal_mac_enable_reg_s_mask : std_logic;
signal internal_mac_subtraction_reg_a_b : std_logic;
signal internal_mac_sel_multiply_two_a_b : std_logic;
signal internal_mac_sel_reg_y_output : std_logic;
signal internal_sm_mac_write_enable_output : std_logic;
signal internal_mac_memory_double_mode : std_logic;
signal internal_mac_memory_only_write_mode : std_logic;
signal internal_base_address_generator_o_increment_previous_address : std_logic;
signal internal_sm_free_flag : std_logic;


-- 0000 multiplication with no reduction
constant first_state_multiplication_direct_operand_size_1 : std_logic_vector(11 downto 0)                                      := std_logic_vector(to_unsigned(0,12));
constant first_state_multiplication_direct_operand_size_2_3_4_5_6_7_8 : std_logic_vector(11 downto 0)                          := std_logic_vector(to_unsigned(2,12));
-- 0001 square with no reduction                                                                                               
constant first_state_square_direct_operand_size_1 : std_logic_vector(11 downto 0)                                              := std_logic_vector(to_unsigned(141,12));
constant first_state_square_direct_operand_size_2_3_4_5_6_7_8 : std_logic_vector(11 downto 0)                                  := std_logic_vector(to_unsigned(143,12));
-- 0010 multiplication with reduction and prime line not equal to 1                                                            
constant first_state_multiplication_with_reduction_operand_size_1 : std_logic_vector(11 downto 0)                              := std_logic_vector(to_unsigned(226,12));
constant first_state_multiplication_with_reduction_operand_size_2_3_4_5_6_7_8 : std_logic_vector(11 downto 0)                  := std_logic_vector(to_unsigned(231,12));
-- 0010 multiplication with reduction and prime line equal to 1                                                     
constant first_state_multiplication_with_reduction_special_prime_1_operand_size_1 : std_logic_vector(11 downto 0)              := std_logic_vector(to_unsigned(510,12));
constant first_state_multiplication_with_reduction_special_prime_1_operand_size_2_3_4_5_6_7_8 : std_logic_vector(11 downto 0)  := std_logic_vector(to_unsigned(513,12));
constant first_state_multiplication_with_reduction_special_prime_2_operand_size_2_3_4_5_6_7_8 : std_logic_vector(11 downto 0)  := std_logic_vector(to_unsigned(765,12));
constant first_state_multiplication_with_reduction_special_prime_3_operand_size_3_4_5_6_7_8 : std_logic_vector(11 downto 0)    := std_logic_vector(to_unsigned(1002,12));
-- 0011 square with reduction and prime line not equal to 1                                                                    
constant first_state_square_with_reduction_operand_size_1 : std_logic_vector(11 downto 0)                                      := std_logic_vector(to_unsigned(1217,12));
constant first_state_square_with_reduction_operand_size_2_3_4_5_6_7_8 : std_logic_vector(11 downto 0)                          := std_logic_vector(to_unsigned(1222,12));
-- 0011 square with reduction and prime line equal to 1                                                                        
constant first_state_square_with_reduction_special_prime_1_operand_size_1 : std_logic_vector(11 downto 0)                      := std_logic_vector(to_unsigned(1445,12));
constant first_state_square_with_reduction_special_prime_1_operand_size_2_3_4_5_6_7_8 : std_logic_vector(11 downto 0)          := std_logic_vector(to_unsigned(1448,12));
constant first_state_square_with_reduction_special_prime_2_operand_size_2_3_4_5_6_7_8 : std_logic_vector(11 downto 0)          := std_logic_vector(to_unsigned(1643,12));
constant first_state_square_with_reduction_special_prime_3_operand_size_3_4_5_6_7_8 : std_logic_vector(11 downto 0)            := std_logic_vector(to_unsigned(1824,12));
-- 0100 addition with no reduction                                                                                             
constant first_state_addition_subtraction_direct_operand_size_1 : std_logic_vector(11 downto 0)                                := std_logic_vector(to_unsigned(1984, 12));
constant first_state_addition_subtraction_direct_operand_size_2_3_4_5_6_7_8 : std_logic_vector(11 downto 0)                    := std_logic_vector(to_unsigned(1986, 12));
-- 0101 iterative modular reduction                                                                                            
constant first_state_iterative_modular_reduction_operand_size_1 : std_logic_vector(11 downto 0)                                := std_logic_vector(to_unsigned(2007, 12));
constant first_state_iterative_modular_reduction_operand_size_2 : std_logic_vector(11 downto 0)                                := std_logic_vector(to_unsigned(2012, 12));
constant first_state_iterative_modular_reduction_operand_size_3 : std_logic_vector(11 downto 0)                                := std_logic_vector(to_unsigned(2020, 12));
constant first_state_iterative_modular_reduction_operand_size_4 : std_logic_vector(11 downto 0)                                := std_logic_vector(to_unsigned(2031, 12));
constant first_state_iterative_modular_reduction_operand_size_5 : std_logic_vector(11 downto 0)                                := std_logic_vector(to_unsigned(2045, 12));
constant first_state_iterative_modular_reduction_operand_size_6 : std_logic_vector(11 downto 0)                                := std_logic_vector(to_unsigned(2062, 12));
constant first_state_iterative_modular_reduction_operand_size_7 : std_logic_vector(11 downto 0)                                := std_logic_vector(to_unsigned(2082, 12));
constant first_state_iterative_modular_reduction_operand_size_8 : std_logic_vector(11 downto 0)                                := std_logic_vector(to_unsigned(2105, 12));
-- 0110 addition with no reduction                                                                                             
constant first_state_addition_subtraction_with_reduction_operand_size_1 : std_logic_vector(11 downto 0)                        := std_logic_vector(to_unsigned(2131, 12));
constant first_state_addition_subtraction_with_reduction_operand_size_2_3_4_5_6_7_8 : std_logic_vector(11 downto 0)            := std_logic_vector(to_unsigned(2136, 12));


type state is (reset, decode_instruction, instruction_execution, multiplication_direct_0, multiplication_direct_2, square_direct_0, square_direct_2, multiplication_with_reduction_special_prime_1_0, multiplication_with_reduction_special_prime_1_3, multiplication_with_reduction_special_prime_2_0, multiplication_with_reduction_special_prime_3_0, multiplication_with_reduction_0, multiplication_with_reduction_5, square_with_reduction_special_prime_1_0, square_with_reduction_special_prime_1_3, square_with_reduction_special_prime_2_0, square_with_reduction_special_prime_3_0, square_with_reduction_0, square_with_reduction_5, addition_subtraction_direct_0, addition_subtraction_direct_2, iterative_modular_reduction_0, iterative_modular_reduction_5, iterative_modular_reduction_13, iterative_modular_reduction_24, iterative_modular_reduction_38, iterative_modular_reduction_55, iterative_modular_reduction_75, iterative_modular_reduction_98, addition_subtraction_with_reduction_0, addition_subtraction_with_reduction_5);

signal actual_state, next_state : state;

signal internal_next_sel_output_rom : std_logic;
signal internal_next_update_rom_address : std_logic;
signal internal_next_sel_load_new_rom_address : std_logic;
signal internal_next_sm_rotation_size : std_logic_vector(1 downto 0);
signal internal_next_sm_circular_shift_enable : std_logic;
signal internal_next_sel_address_a : std_logic;
signal internal_next_sel_address_b_prime : std_logic_vector(1 downto 0);
signal internal_next_sm_specific_mac_address_a : std_logic_vector(2 downto 0);
signal internal_next_sm_specific_mac_address_b : std_logic_vector(2 downto 0);
signal internal_next_sm_specific_mac_address_o : std_logic_vector(2 downto 0);
signal internal_next_sm_specific_mac_next_address_o : std_logic_vector(2 downto 0);
signal internal_next_mac_enable_signed_a : std_logic;
signal internal_next_mac_enable_signed_b : std_logic;
signal internal_next_mac_sel_load_reg_a : std_logic_vector(1 downto 0);
signal internal_next_mac_clear_reg_b : std_logic;
signal internal_next_mac_clear_reg_acc : std_logic;
signal internal_next_mac_sel_shift_reg_o : std_logic;
signal internal_next_mac_enable_update_reg_s : std_logic;
signal internal_next_mac_sel_reg_s_reg_o_sign : std_logic;
signal internal_next_mac_reg_s_reg_o_positive : std_logic;
signal internal_next_sm_sign_a_mode : std_logic;
signal internal_next_sm_mac_operation_mode : std_logic_vector(1 downto 0);
signal internal_next_mac_enable_reg_s_mask : std_logic;
signal internal_next_mac_subtraction_reg_a_b : std_logic;
signal internal_next_mac_sel_multiply_two_a_b : std_logic;
signal internal_next_mac_sel_reg_y_output : std_logic;
signal internal_next_sm_mac_write_enable_output : std_logic;
signal internal_next_mac_memory_double_mode : std_logic;
signal internal_next_mac_memory_only_write_mode : std_logic;
signal internal_next_base_address_generator_o_increment_previous_address : std_logic;
signal internal_next_sm_free_flag : std_logic;

signal reg_rom_last_state : std_logic;

begin

registers_state : process(clk, rstn)
begin
    if(rstn = '0') then
        actual_state <= reset;
    elsif(rising_edge(clk)) then
        actual_state <= next_state;
    end if;
end process;

registers_state_output : process(clk)
begin
    if(rising_edge(clk)) then
        if(rstn = '0') then
            internal_sel_output_rom <= '0';
            internal_update_rom_address <= '1';
            internal_sel_load_new_rom_address <= '1';
            internal_sm_rotation_size <= "11";
            internal_sm_circular_shift_enable <= '0';
            internal_sel_address_a <= '0';
            internal_sel_address_b_prime <= "00";
            internal_sm_specific_mac_address_a <= "000";
            internal_sm_specific_mac_address_b <= "000";
            internal_sm_specific_mac_address_o <= "000";
            internal_sm_specific_mac_next_address_o <= "001";
            internal_mac_enable_signed_a <= '0';
            internal_mac_enable_signed_b <= '0';
            internal_mac_sel_load_reg_a <= "00";
            internal_mac_clear_reg_b <= '0';
            internal_mac_clear_reg_acc <= '0';
            internal_mac_sel_shift_reg_o <= '0';
            internal_mac_enable_update_reg_s <= '0';
            internal_mac_sel_reg_s_reg_o_sign <= '0';
            internal_mac_reg_s_reg_o_positive <= '0';
            internal_sm_sign_a_mode <= '0';
            internal_sm_mac_operation_mode <= "00";
            internal_mac_enable_reg_s_mask <= '0';
            internal_mac_subtraction_reg_a_b <= '0';
            internal_mac_sel_multiply_two_a_b <= '0';
            internal_mac_sel_reg_y_output <= '0';
            internal_sm_mac_write_enable_output <= '0';
            internal_mac_memory_double_mode <= '0';
            internal_mac_memory_only_write_mode <= '0';
            internal_base_address_generator_o_increment_previous_address <= '0';
            internal_sm_free_flag <= '0';
        else
            internal_sel_output_rom <= internal_next_sel_output_rom;
            internal_update_rom_address <= internal_next_update_rom_address;
            internal_sel_load_new_rom_address <= internal_next_sel_load_new_rom_address;
            if(internal_sel_output_rom = '1') then
                internal_sm_rotation_size <= rom_sm_rotation_size;
                internal_sm_circular_shift_enable <= internal_next_sm_circular_shift_enable;
                internal_sel_address_a <= rom_sel_address_a;
                internal_sel_address_b_prime <= rom_sel_address_b_prime;
                internal_sm_specific_mac_address_a <= rom_sm_specific_mac_address_a;
                internal_sm_specific_mac_address_b <= rom_sm_specific_mac_address_b;
                internal_sm_specific_mac_address_o <= rom_sm_specific_mac_address_o;
                internal_sm_specific_mac_next_address_o <= rom_sm_specific_mac_next_address_o;
                internal_mac_enable_signed_a <= rom_mac_enable_signed_a;
                internal_mac_enable_signed_b <= rom_mac_enable_signed_b;
                internal_mac_sel_load_reg_a <= rom_mac_sel_load_reg_a;
                internal_mac_clear_reg_b <= rom_mac_clear_reg_b;
                internal_mac_clear_reg_acc <= rom_mac_clear_reg_acc;
                internal_mac_sel_shift_reg_o <= rom_mac_sel_shift_reg_o;
                internal_mac_enable_update_reg_s <= rom_mac_enable_update_reg_s;
                internal_mac_sel_reg_s_reg_o_sign <= rom_mac_sel_reg_s_reg_o_sign;
                internal_mac_reg_s_reg_o_positive <= rom_mac_reg_s_reg_o_positive;
                internal_sm_sign_a_mode <= rom_sm_sign_a_mode;
                internal_sm_mac_operation_mode <= rom_sm_mac_operation_mode;
                internal_mac_enable_reg_s_mask <= rom_mac_enable_reg_s_mask;
                internal_mac_subtraction_reg_a_b <= rom_mac_subtraction_reg_a_b;
                internal_mac_sel_multiply_two_a_b <= rom_mac_sel_multiply_two_a_b;
                internal_mac_sel_reg_y_output <= rom_mac_sel_reg_y_output;
                internal_sm_mac_write_enable_output <= rom_sm_mac_write_enable_output;
                internal_mac_memory_double_mode <= rom_mac_memory_double_mode;
                internal_mac_memory_only_write_mode <= rom_mac_memory_only_write_mode;
                internal_base_address_generator_o_increment_previous_address <= rom_base_address_generator_o_increment_previous_address;
                internal_sm_free_flag <= internal_next_sm_free_flag;
            else
                internal_sm_rotation_size <= internal_next_sm_rotation_size;
                internal_sm_circular_shift_enable <= internal_next_sm_circular_shift_enable;
                internal_sel_address_a <= internal_next_sel_address_a;
                internal_sel_address_b_prime <= internal_next_sel_address_b_prime;
                internal_sm_specific_mac_address_a <= internal_next_sm_specific_mac_address_a;
                internal_sm_specific_mac_address_b <= internal_next_sm_specific_mac_address_b;
                internal_sm_specific_mac_address_o <= internal_next_sm_specific_mac_address_o;
                internal_sm_specific_mac_next_address_o <= internal_next_sm_specific_mac_next_address_o;
                internal_mac_enable_signed_a <= internal_next_mac_enable_signed_a;
                internal_mac_enable_signed_b <= internal_next_mac_enable_signed_b;
                internal_mac_sel_load_reg_a <= internal_next_mac_sel_load_reg_a;
                internal_mac_clear_reg_b <= internal_next_mac_clear_reg_b;
                internal_mac_clear_reg_acc <= internal_next_mac_clear_reg_acc;
                internal_mac_sel_shift_reg_o <= internal_next_mac_sel_shift_reg_o;
                internal_mac_enable_update_reg_s <= internal_next_mac_enable_update_reg_s;
                internal_mac_sel_reg_s_reg_o_sign <= internal_next_mac_sel_reg_s_reg_o_sign;
                internal_mac_reg_s_reg_o_positive <= internal_next_mac_reg_s_reg_o_positive;
                internal_sm_sign_a_mode <= internal_next_sm_sign_a_mode;
                internal_sm_mac_operation_mode <= internal_next_sm_mac_operation_mode;
                internal_mac_enable_reg_s_mask <= internal_next_mac_enable_reg_s_mask;
                internal_mac_subtraction_reg_a_b <= internal_next_mac_subtraction_reg_a_b;
                internal_mac_sel_multiply_two_a_b <= internal_next_mac_sel_multiply_two_a_b;
                internal_mac_sel_reg_y_output <= internal_next_mac_sel_reg_y_output;
                internal_sm_mac_write_enable_output <= internal_next_sm_mac_write_enable_output;
                internal_mac_memory_double_mode <= internal_next_mac_memory_double_mode;
                internal_mac_memory_only_write_mode <= internal_next_mac_memory_only_write_mode;
                internal_base_address_generator_o_increment_previous_address <= internal_next_base_address_generator_o_increment_previous_address;
                internal_sm_free_flag <= internal_next_sm_free_flag;
            end if;
        end if;
    end if;
end process;

update_output : process(next_state)
begin
    case (next_state) is
        when reset =>
            internal_next_sel_output_rom <= '0';
            internal_next_update_rom_address <= '1';
            internal_next_sel_load_new_rom_address <= '1';
            internal_next_sm_rotation_size <= "11";
            internal_next_sm_circular_shift_enable <= '0';
            internal_next_sel_address_a <= '0';
            internal_next_sel_address_b_prime <= "00";
            internal_next_sm_specific_mac_address_a <= "000";
            internal_next_sm_specific_mac_address_b <= "000";
            internal_next_sm_specific_mac_address_o <= "000";
            internal_next_sm_specific_mac_next_address_o <= "001";
            internal_next_mac_enable_signed_a <= '0';
            internal_next_mac_enable_signed_b <= '0';
            internal_next_mac_sel_load_reg_a <= "11";
            internal_next_mac_clear_reg_b <= '1';
            internal_next_mac_clear_reg_acc <= '1';
            internal_next_mac_sel_shift_reg_o <= '0';
            internal_next_mac_enable_update_reg_s <= '0';
            internal_next_mac_sel_reg_s_reg_o_sign <= '0';
            internal_next_mac_reg_s_reg_o_positive <= '0';
            internal_next_sm_sign_a_mode <= '0';
            internal_next_sm_mac_operation_mode <= "10";
            internal_next_mac_enable_reg_s_mask <= '0';
            internal_next_mac_subtraction_reg_a_b <= '0';
            internal_next_mac_sel_multiply_two_a_b <= '0';
            internal_next_mac_sel_reg_y_output <= '0';
            internal_next_sm_mac_write_enable_output <= '0';
            internal_next_mac_memory_double_mode <= '0';
            internal_next_mac_memory_only_write_mode <= '0';
            internal_next_base_address_generator_o_increment_previous_address <= '0';
            internal_next_sm_free_flag <= '1';
        when decode_instruction =>
            internal_next_sel_output_rom <= '0';
            internal_next_update_rom_address <= '1';
            internal_next_sel_load_new_rom_address <= '1';
            internal_next_sm_free_flag <= '1';
            internal_next_sm_rotation_size <= "11";
            internal_next_sm_circular_shift_enable <= '0';
            internal_next_sel_address_a <= '0';
            internal_next_sel_address_b_prime <= "00";
            internal_next_sm_specific_mac_address_a <= "000";
            internal_next_sm_specific_mac_address_b <= "000";
            internal_next_sm_specific_mac_address_o <= "000";
            internal_next_sm_specific_mac_next_address_o <= "001";
            internal_next_mac_enable_signed_a <= '0';
            internal_next_mac_enable_signed_b <= '0';
            internal_next_mac_sel_load_reg_a <= "11";
            internal_next_mac_clear_reg_b <= '1';
            internal_next_mac_clear_reg_acc <= '1';
            internal_next_mac_sel_shift_reg_o <= '0';
            internal_next_mac_enable_update_reg_s <= '0';
            internal_next_mac_sel_reg_s_reg_o_sign <= '0';
            internal_next_mac_reg_s_reg_o_positive <= '0';
            internal_next_sm_sign_a_mode <= '0';
            internal_next_sm_mac_operation_mode <= "10";
            internal_next_mac_enable_reg_s_mask <= '0';
            internal_next_mac_subtraction_reg_a_b <= '0';
            internal_next_mac_sel_multiply_two_a_b <= '0';
            internal_next_mac_sel_reg_y_output <= '0';
            internal_next_sm_mac_write_enable_output <= '0';
            internal_next_mac_memory_double_mode <= '0';
            internal_next_mac_memory_only_write_mode <= '0';
            internal_next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_0 =>
            -- -- In case of size 1
            -- reg_a = a0_X; reg_b = b0_X; reg_acc = 0; o0_X = reg_o; o1_X = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
            internal_next_sel_output_rom <= '1';
            internal_next_update_rom_address <= '1';
            internal_next_sel_load_new_rom_address <= '0';
            internal_next_sm_free_flag <= '0';
            internal_next_sm_rotation_size <= "11";
            internal_next_sm_circular_shift_enable <= '1';
            internal_next_sel_address_a <= '0';
            internal_next_sel_address_b_prime <= "00";
            internal_next_sm_specific_mac_address_a <= "000";
            internal_next_sm_specific_mac_address_b <= "000";
            internal_next_sm_specific_mac_address_o <= "000";
            internal_next_sm_specific_mac_next_address_o <= "001";
            internal_next_mac_enable_signed_a <= '1';
            internal_next_mac_enable_signed_b <= '1';
            internal_next_mac_sel_load_reg_a <= "00";
            internal_next_mac_clear_reg_b <= '0';
            internal_next_mac_clear_reg_acc <= '1';
            internal_next_mac_sel_shift_reg_o <= '0';
            internal_next_mac_enable_update_reg_s <= '0';
            internal_next_mac_sel_reg_s_reg_o_sign <= '0';
            internal_next_mac_reg_s_reg_o_positive <= '0';
            internal_next_sm_sign_a_mode <= '0';
            internal_next_sm_mac_operation_mode <= "10";
            internal_next_mac_enable_reg_s_mask <= '0';
            internal_next_mac_subtraction_reg_a_b <= '0';
            internal_next_mac_sel_multiply_two_a_b <= '0';
            internal_next_mac_sel_reg_y_output <= '0';
            internal_next_sm_mac_write_enable_output <= '1';
            internal_next_mac_memory_double_mode <= '1';
            internal_next_mac_memory_only_write_mode <= '1';
            internal_next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_2 =>
            -- -- Other cases
            -- reg_a = a0_X; reg_b = b0_X; reg_acc = 0; o0_X = reg_o; operation : a*b + acc; o0_X = reg_o;
            internal_next_sel_output_rom <= '1';
            internal_next_update_rom_address <= '1';
            internal_next_sel_load_new_rom_address <= '0';
            internal_next_sm_free_flag <= '0';
            internal_next_sm_rotation_size <= "11";
            internal_next_sm_circular_shift_enable <= '1';
            internal_next_sel_address_a <= '0';
            internal_next_sel_address_b_prime <= "00";
            internal_next_sm_specific_mac_address_a <= "000";
            internal_next_sm_specific_mac_address_b <= "000";
            internal_next_sm_specific_mac_address_o <= "000";
            internal_next_sm_specific_mac_next_address_o <= "001";
            internal_next_mac_enable_signed_a <= '0';
            internal_next_mac_enable_signed_b <= '0';
            internal_next_mac_sel_load_reg_a <= "00";
            internal_next_mac_clear_reg_b <= '0';
            internal_next_mac_clear_reg_acc <= '1';
            internal_next_mac_sel_shift_reg_o <= '0';
            internal_next_mac_enable_update_reg_s <= '0';
            internal_next_mac_sel_reg_s_reg_o_sign <= '0';
            internal_next_mac_reg_s_reg_o_positive <= '0';
            internal_next_sm_sign_a_mode <= '0';
            internal_next_sm_mac_operation_mode <= "10";
            internal_next_mac_enable_reg_s_mask <= '0';
            internal_next_mac_subtraction_reg_a_b <= '0';
            internal_next_mac_sel_multiply_two_a_b <= '0';
            internal_next_mac_sel_reg_y_output <= '0';
            internal_next_sm_mac_write_enable_output <= '1';
            internal_next_mac_memory_double_mode <= '0';
            internal_next_mac_memory_only_write_mode <= '0';
            internal_next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_0 => 
            -- -- In case of size 1
            -- reg_a = a0_X; reg_b = a0_X; reg_acc = 0; o0_X = reg_o; o1_X = reg_o >> 256; Enable sign a,b; operation : a*b + acc;
            internal_next_sel_output_rom <= '1';
            internal_next_update_rom_address <= '1';
            internal_next_sel_load_new_rom_address <= '0';
            internal_next_sm_free_flag <= '0';
            internal_next_sm_rotation_size <= "11";
            internal_next_sm_circular_shift_enable <= '1';
            internal_next_sel_address_a <= '0';
            internal_next_sel_address_b_prime <= "00";
            internal_next_sm_specific_mac_address_a <= "000";
            internal_next_sm_specific_mac_address_b <= "000";
            internal_next_sm_specific_mac_address_o <= "000";
            internal_next_sm_specific_mac_next_address_o <= "001";
            internal_next_mac_enable_signed_a <= '1';
            internal_next_mac_enable_signed_b <= '1';
            internal_next_mac_sel_load_reg_a <= "00";
            internal_next_mac_clear_reg_b <= '0';
            internal_next_mac_clear_reg_acc <= '1';
            internal_next_mac_sel_shift_reg_o <= '0';
            internal_next_mac_enable_update_reg_s <= '0';
            internal_next_mac_sel_reg_s_reg_o_sign <= '0';
            internal_next_mac_reg_s_reg_o_positive <= '0';
            internal_next_sm_sign_a_mode <= '0';
            internal_next_sm_mac_operation_mode <= "10";
            internal_next_mac_enable_reg_s_mask <= '0';
            internal_next_mac_subtraction_reg_a_b <= '0';
            internal_next_mac_sel_multiply_two_a_b <= '0';
            internal_next_mac_sel_reg_y_output <= '0';
            internal_next_sm_mac_write_enable_output <= '1';
            internal_next_mac_memory_double_mode <= '1';
            internal_next_mac_memory_only_write_mode <= '1';
            internal_next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_2 => 
            -- -- In case of sizes 2, 3, 4, 5, 6, 7, 8
            -- reg_a = a0_X; reg_b = a0_X; reg_acc = 0; o0_X = reg_o; operation : a*b + acc;
            internal_next_sel_output_rom <= '1';
            internal_next_update_rom_address <= '1';
            internal_next_sel_load_new_rom_address <= '0';
            internal_next_sm_free_flag <= '0';
            internal_next_sm_rotation_size <= "11";
            internal_next_sm_circular_shift_enable <= '1';
            internal_next_sel_address_a <= '0';
            internal_next_sel_address_b_prime <= "00";
            internal_next_sm_specific_mac_address_a <= "000";
            internal_next_sm_specific_mac_address_b <= "000";
            internal_next_sm_specific_mac_address_o <= "000";
            internal_next_sm_specific_mac_next_address_o <= "001";
            internal_next_mac_enable_signed_a <= '0';
            internal_next_mac_enable_signed_b <= '0';
            internal_next_mac_sel_load_reg_a <= "00";
            internal_next_mac_clear_reg_b <= '0';
            internal_next_mac_clear_reg_acc <= '1';
            internal_next_mac_sel_shift_reg_o <= '0';
            internal_next_mac_enable_update_reg_s <= '0';
            internal_next_mac_sel_reg_s_reg_o_sign <= '0';
            internal_next_mac_reg_s_reg_o_positive <= '0';
            internal_next_sm_sign_a_mode <= '0';
            internal_next_sm_mac_operation_mode <= "10";
            internal_next_mac_enable_reg_s_mask <= '0';
            internal_next_mac_subtraction_reg_a_b <= '0';
            internal_next_mac_sel_multiply_two_a_b <= '0';
            internal_next_mac_sel_reg_y_output <= '0';
            internal_next_sm_mac_write_enable_output <= '1';
            internal_next_mac_memory_double_mode <= '0';
            internal_next_mac_memory_only_write_mode <= '0';
            internal_next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_0 =>
            -- -- In case of size 1
            -- reg_a = a0_X; reg_b = b0_X; reg_acc = 0; Enable sign a,b; operation : a*b + acc;
            internal_next_sel_output_rom <= '1';
            internal_next_update_rom_address <= '1';
            internal_next_sel_load_new_rom_address <= '0';
            internal_next_sm_free_flag <= '0';
            internal_next_sm_rotation_size <= "11";
            internal_next_sm_circular_shift_enable <= '1';
            internal_next_sel_address_a <= '0';
            internal_next_sel_address_b_prime <= "00";
            internal_next_sm_specific_mac_address_a <= "000";
            internal_next_sm_specific_mac_address_b <= "000";
            internal_next_sm_specific_mac_address_o <= "000";
            internal_next_sm_specific_mac_next_address_o <= "001";
            internal_next_mac_enable_signed_a <= '0';
            internal_next_mac_enable_signed_b <= '0';
            internal_next_mac_sel_load_reg_a <= "00";
            internal_next_mac_clear_reg_b <= '0';
            internal_next_mac_clear_reg_acc <= '1';
            internal_next_mac_sel_shift_reg_o <= '0';
            internal_next_mac_enable_update_reg_s <= '0';
            internal_next_mac_sel_reg_s_reg_o_sign <= '0';
            internal_next_mac_reg_s_reg_o_positive <= '0';
            internal_next_sm_sign_a_mode <= '0';
            internal_next_sm_mac_operation_mode <= "10";
            internal_next_mac_enable_reg_s_mask <= '0';
            internal_next_mac_subtraction_reg_a_b <= '0';
            internal_next_mac_sel_multiply_two_a_b <= '0';
            internal_next_mac_sel_reg_y_output <= '0';
            internal_next_sm_mac_write_enable_output <= '0';
            internal_next_mac_memory_double_mode <= '0';
            internal_next_mac_memory_only_write_mode <= '0';
            internal_next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1_3 =>
            -- -- In case of sizes 2, 3, 4, 5, 6, 7, 8
            -- reg_a = a0_X; reg_b = b0_X; reg_acc = 0; o0_X = reg_o; operation : a*b + acc;
            internal_next_sel_output_rom <= '1';
            internal_next_update_rom_address <= '1';
            internal_next_sel_load_new_rom_address <= '0';
            internal_next_sm_free_flag <= '0';
            internal_next_sm_rotation_size <= "11";
            internal_next_sm_circular_shift_enable <= '1';
            internal_next_sel_address_a <= '0';
            internal_next_sel_address_b_prime <= "00";
            internal_next_sm_specific_mac_address_a <= "000";
            internal_next_sm_specific_mac_address_b <= "000";
            internal_next_sm_specific_mac_address_o <= "000";
            internal_next_sm_specific_mac_next_address_o <= "001";
            internal_next_mac_enable_signed_a <= '0';
            internal_next_mac_enable_signed_b <= '0';
            internal_next_mac_sel_load_reg_a <= "00";
            internal_next_mac_clear_reg_b <= '0';
            internal_next_mac_clear_reg_acc <= '1';
            internal_next_mac_sel_shift_reg_o <= '0';
            internal_next_mac_enable_update_reg_s <= '0';
            internal_next_mac_sel_reg_s_reg_o_sign <= '0';
            internal_next_mac_reg_s_reg_o_positive <= '0';
            internal_next_sm_sign_a_mode <= '0';
            internal_next_sm_mac_operation_mode <= "10";
            internal_next_mac_enable_reg_s_mask <= '0';
            internal_next_mac_subtraction_reg_a_b <= '0';
            internal_next_mac_sel_multiply_two_a_b <= '0';
            internal_next_mac_sel_reg_y_output <= '0';
            internal_next_sm_mac_write_enable_output <= '1';
            internal_next_mac_memory_double_mode <= '0';
            internal_next_mac_memory_only_write_mode <= '0';
            internal_next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_2_0 =>
            -- With 2 zeroes in prime sharp
            -- -- In case of sizes 2, 3, 4, 5, 6, 7, 8
            -- reg_a = a0_X; reg_b = b0_X; reg_acc = 0; o0_X = reg_o; operation : a*b + acc;
            internal_next_sel_output_rom <= '1';
            internal_next_update_rom_address <= '1';
            internal_next_sel_load_new_rom_address <= '0';
            internal_next_sm_free_flag <= '0';
            internal_next_sm_rotation_size <= "11";
            internal_next_sm_circular_shift_enable <= '1';
            internal_next_sel_address_a <= '0';
            internal_next_sel_address_b_prime <= "00";
            internal_next_sm_specific_mac_address_a <= "000";
            internal_next_sm_specific_mac_address_b <= "000";
            internal_next_sm_specific_mac_address_o <= "000";
            internal_next_sm_specific_mac_next_address_o <= "001";
            internal_next_mac_enable_signed_a <= '0';
            internal_next_mac_enable_signed_b <= '0';
            internal_next_mac_sel_load_reg_a <= "00";
            internal_next_mac_clear_reg_b <= '0';
            internal_next_mac_clear_reg_acc <= '1';
            internal_next_mac_sel_shift_reg_o <= '0';
            internal_next_mac_enable_update_reg_s <= '0';
            internal_next_mac_sel_reg_s_reg_o_sign <= '0';
            internal_next_mac_reg_s_reg_o_positive <= '0';
            internal_next_sm_sign_a_mode <= '0';
            internal_next_sm_mac_operation_mode <= "10";
            internal_next_mac_enable_reg_s_mask <= '0';
            internal_next_mac_subtraction_reg_a_b <= '0';
            internal_next_mac_sel_multiply_two_a_b <= '0';
            internal_next_mac_sel_reg_y_output <= '0';
            internal_next_sm_mac_write_enable_output <= '1';
            internal_next_mac_memory_double_mode <= '0';
            internal_next_mac_memory_only_write_mode <= '0';
            internal_next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3_0 =>
            -- -- In case of sizes 3, 4, 5, 6, 7, 8
            -- reg_a = a0_X; reg_b = b0_X; reg_acc = 0; o0_X = reg_o; operation : a*b + acc;
            internal_next_sel_output_rom <= '1';
            internal_next_update_rom_address <= '1';
            internal_next_sel_load_new_rom_address <= '0';
            internal_next_sm_free_flag <= '0';
            internal_next_sm_rotation_size <= "11";
            internal_next_sm_circular_shift_enable <= '1';
            internal_next_sel_address_a <= '0';
            internal_next_sel_address_b_prime <= "00";
            internal_next_sm_specific_mac_address_a <= "000";
            internal_next_sm_specific_mac_address_b <= "000";
            internal_next_sm_specific_mac_address_o <= "000";
            internal_next_sm_specific_mac_next_address_o <= "001";
            internal_next_mac_enable_signed_a <= '0';
            internal_next_mac_enable_signed_b <= '0';
            internal_next_mac_sel_load_reg_a <= "00";
            internal_next_mac_clear_reg_b <= '0';
            internal_next_mac_clear_reg_acc <= '1';
            internal_next_mac_sel_shift_reg_o <= '0';
            internal_next_mac_enable_update_reg_s <= '0';
            internal_next_mac_sel_reg_s_reg_o_sign <= '0';
            internal_next_mac_reg_s_reg_o_positive <= '0';
            internal_next_sm_sign_a_mode <= '0';
            internal_next_sm_mac_operation_mode <= "10";
            internal_next_mac_enable_reg_s_mask <= '0';
            internal_next_mac_subtraction_reg_a_b <= '0';
            internal_next_mac_sel_multiply_two_a_b <= '0';
            internal_next_mac_sel_reg_y_output <= '0';
            internal_next_sm_mac_write_enable_output <= '1';
            internal_next_mac_memory_double_mode <= '0';
            internal_next_mac_memory_only_write_mode <= '0';
            internal_next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_0 =>
            -- -- In case of size 1
            -- reg_a = a0_X; reg_b = b0_X; reg_acc = 0; Enable sign a,b; operation : a*b + acc;
            internal_next_sel_output_rom <= '1';
            internal_next_update_rom_address <= '1';
            internal_next_sel_load_new_rom_address <= '0';
            internal_next_sm_free_flag <= '0';
            internal_next_sm_rotation_size <= "11";
            internal_next_sm_circular_shift_enable <= '1';
            internal_next_sel_address_a <= '0';
            internal_next_sel_address_b_prime <= "00";
            internal_next_sm_specific_mac_address_a <= "000";
            internal_next_sm_specific_mac_address_b <= "000";
            internal_next_sm_specific_mac_address_o <= "000";
            internal_next_sm_specific_mac_next_address_o <= "001";
            internal_next_mac_enable_signed_a <= '1';
            internal_next_mac_enable_signed_b <= '1';
            internal_next_mac_sel_load_reg_a <= "00";
            internal_next_mac_clear_reg_b <= '0';
            internal_next_mac_clear_reg_acc <= '1';
            internal_next_mac_sel_shift_reg_o <= '0';
            internal_next_mac_enable_update_reg_s <= '0';
            internal_next_mac_sel_reg_s_reg_o_sign <= '0';
            internal_next_mac_reg_s_reg_o_positive <= '0';
            internal_next_sm_sign_a_mode <= '0';
            internal_next_sm_mac_operation_mode <= "10";
            internal_next_mac_enable_reg_s_mask <= '0';
            internal_next_mac_subtraction_reg_a_b <= '0';
            internal_next_mac_sel_multiply_two_a_b <= '0';
            internal_next_mac_sel_reg_y_output <= '0';
            internal_next_sm_mac_write_enable_output <= '0';
            internal_next_mac_memory_double_mode <= '0';
            internal_next_mac_memory_only_write_mode <= '0';
            internal_next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_5 =>
            -- -- In case of sizes 2, 3, 4, 5, 6, 7, 8
            -- reg_a = a0_X; reg_b = b0_X; reg_acc = 0; operation : a*b + acc;
            internal_next_sel_output_rom <= '1';
            internal_next_update_rom_address <= '1';
            internal_next_sel_load_new_rom_address <= '0';
            internal_next_sm_free_flag <= '0';
            internal_next_sm_rotation_size <= "11";
            internal_next_sm_circular_shift_enable <= '1';
            internal_next_sel_address_a <= '0';
            internal_next_sel_address_b_prime <= "00";
            internal_next_sm_specific_mac_address_a <= "000";
            internal_next_sm_specific_mac_address_b <= "000";
            internal_next_sm_specific_mac_address_o <= "000";
            internal_next_sm_specific_mac_next_address_o <= "001";
            internal_next_mac_enable_signed_a <= '0';
            internal_next_mac_enable_signed_b <= '0';
            internal_next_mac_sel_load_reg_a <= "00";
            internal_next_mac_clear_reg_b <= '0';
            internal_next_mac_clear_reg_acc <= '1';
            internal_next_mac_sel_shift_reg_o <= '0';
            internal_next_mac_enable_update_reg_s <= '0';
            internal_next_mac_sel_reg_s_reg_o_sign <= '0';
            internal_next_mac_reg_s_reg_o_positive <= '0';
            internal_next_sm_sign_a_mode <= '0';
            internal_next_sm_mac_operation_mode <= "10";
            internal_next_mac_enable_reg_s_mask <= '0';
            internal_next_mac_subtraction_reg_a_b <= '0';
            internal_next_mac_sel_multiply_two_a_b <= '0';
            internal_next_mac_sel_reg_y_output <= '0';
            internal_next_sm_mac_write_enable_output <= '0';
            internal_next_mac_memory_double_mode <= '0';
            internal_next_mac_memory_only_write_mode <= '0';
            internal_next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_0 =>
            -- -- In case of size 1
            -- reg_a = a0_X; reg_b = a0_X; reg_acc = 0; Enable sign a,b; operation : a*b + acc;
            internal_next_sel_output_rom <= '1';
            internal_next_update_rom_address <= '1';
            internal_next_sel_load_new_rom_address <= '0';
            internal_next_sm_free_flag <= '0';
            internal_next_sm_rotation_size <= "11";
            internal_next_sm_circular_shift_enable <= '1';
            internal_next_sel_address_a <= '0';
            internal_next_sel_address_b_prime <= "00";
            internal_next_sm_specific_mac_address_a <= "000";
            internal_next_sm_specific_mac_address_b <= "000";
            internal_next_sm_specific_mac_address_o <= "000";
            internal_next_sm_specific_mac_next_address_o <= "001";
            internal_next_mac_enable_signed_a <= '1';
            internal_next_mac_enable_signed_b <= '1';
            internal_next_mac_sel_load_reg_a <= "00";
            internal_next_mac_clear_reg_b <= '0';
            internal_next_mac_clear_reg_acc <= '1';
            internal_next_mac_sel_shift_reg_o <= '0';
            internal_next_mac_enable_update_reg_s <= '0';
            internal_next_mac_sel_reg_s_reg_o_sign <= '0';
            internal_next_mac_reg_s_reg_o_positive <= '0';
            internal_next_sm_sign_a_mode <= '0';
            internal_next_sm_mac_operation_mode <= "10";
            internal_next_mac_enable_reg_s_mask <= '0';
            internal_next_mac_subtraction_reg_a_b <= '0';
            internal_next_mac_sel_multiply_two_a_b <= '0';
            internal_next_mac_sel_reg_y_output <= '0';
            internal_next_sm_mac_write_enable_output <= '0';
            internal_next_mac_memory_double_mode <= '0';
            internal_next_mac_memory_only_write_mode <= '0';
            internal_next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1_3 =>
            -- -- In case of size 2, 3, 4
            -- reg_a = a0_X; reg_b = a0_X; reg_acc = 0; o0_X = reg_o; operation : a*b + acc;
            internal_next_sel_output_rom <= '1';
            internal_next_update_rom_address <= '1';
            internal_next_sel_load_new_rom_address <= '0';
            internal_next_sm_free_flag <= '0';
            internal_next_sm_rotation_size <= "11";
            internal_next_sm_circular_shift_enable <= '1';
            internal_next_sel_address_a <= '0';
            internal_next_sel_address_b_prime <= "00";
            internal_next_sm_specific_mac_address_a <= "000";
            internal_next_sm_specific_mac_address_b <= "000";
            internal_next_sm_specific_mac_address_o <= "000";
            internal_next_sm_specific_mac_next_address_o <= "001";
            internal_next_mac_enable_signed_a <= '0';
            internal_next_mac_enable_signed_b <= '0';
            internal_next_mac_sel_load_reg_a <= "00";
            internal_next_mac_clear_reg_b <= '0';
            internal_next_mac_clear_reg_acc <= '1';
            internal_next_mac_sel_shift_reg_o <= '0';
            internal_next_mac_enable_update_reg_s <= '0';
            internal_next_mac_sel_reg_s_reg_o_sign <= '0';
            internal_next_mac_reg_s_reg_o_positive <= '0';
            internal_next_sm_sign_a_mode <= '0';
            internal_next_sm_mac_operation_mode <= "10";
            internal_next_mac_enable_reg_s_mask <= '0';
            internal_next_mac_subtraction_reg_a_b <= '0';
            internal_next_mac_sel_multiply_two_a_b <= '0';
            internal_next_mac_sel_reg_y_output <= '0';
            internal_next_sm_mac_write_enable_output <= '1';
            internal_next_mac_memory_double_mode <= '0';
            internal_next_mac_memory_only_write_mode <= '0';
            internal_next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_2_0 =>
            -- -- In case of size 2, 3, 4, 5, 6, 7, 8
            -- reg_a = a0_X; reg_b = a0_X; reg_acc = 0; o0_X = reg_o; operation : a*b + acc;
            internal_next_sel_output_rom <= '1';
            internal_next_update_rom_address <= '1';
            internal_next_sel_load_new_rom_address <= '0';
            internal_next_sm_free_flag <= '0';
            internal_next_sm_rotation_size <= "11";
            internal_next_sm_circular_shift_enable <= '1';
            internal_next_sel_address_a <= '0';
            internal_next_sel_address_b_prime <= "00";
            internal_next_sm_specific_mac_address_a <= "000";
            internal_next_sm_specific_mac_address_b <= "000";
            internal_next_sm_specific_mac_address_o <= "000";
            internal_next_sm_specific_mac_next_address_o <= "001";
            internal_next_mac_enable_signed_a <= '0';
            internal_next_mac_enable_signed_b <= '0';
            internal_next_mac_sel_load_reg_a <= "00";
            internal_next_mac_clear_reg_b <= '0';
            internal_next_mac_clear_reg_acc <= '1';
            internal_next_mac_sel_shift_reg_o <= '0';
            internal_next_mac_enable_update_reg_s <= '0';
            internal_next_mac_sel_reg_s_reg_o_sign <= '0';
            internal_next_mac_reg_s_reg_o_positive <= '0';
            internal_next_sm_sign_a_mode <= '0';
            internal_next_sm_mac_operation_mode <= "10";
            internal_next_mac_enable_reg_s_mask <= '0';
            internal_next_mac_subtraction_reg_a_b <= '0';
            internal_next_mac_sel_multiply_two_a_b <= '0';
            internal_next_mac_sel_reg_y_output <= '0';
            internal_next_sm_mac_write_enable_output <= '1';
            internal_next_mac_memory_double_mode <= '0';
            internal_next_mac_memory_only_write_mode <= '0';
            internal_next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3_0 =>
            -- -- In case of sizes 3, 4, 5, 6, 7, 8
            -- reg_a = a0_X; reg_b = a0_X; reg_acc = 0; o0_X = reg_o; operation : a*b + acc;
            internal_next_sel_output_rom <= '1';
            internal_next_update_rom_address <= '1';
            internal_next_sel_load_new_rom_address <= '0';
            internal_next_sm_free_flag <= '0';
            internal_next_sm_rotation_size <= "11";
            internal_next_sm_circular_shift_enable <= '1';
            internal_next_sel_address_a <= '0';
            internal_next_sel_address_b_prime <= "00";
            internal_next_sm_specific_mac_address_a <= "000";
            internal_next_sm_specific_mac_address_b <= "000";
            internal_next_sm_specific_mac_address_o <= "000";
            internal_next_sm_specific_mac_next_address_o <= "001";
            internal_next_mac_enable_signed_a <= '0';
            internal_next_mac_enable_signed_b <= '0';
            internal_next_mac_sel_load_reg_a <= "00";
            internal_next_mac_clear_reg_b <= '0';
            internal_next_mac_clear_reg_acc <= '1';
            internal_next_mac_sel_shift_reg_o <= '0';
            internal_next_mac_enable_update_reg_s <= '0';
            internal_next_mac_sel_reg_s_reg_o_sign <= '0';
            internal_next_mac_reg_s_reg_o_positive <= '0';
            internal_next_sm_sign_a_mode <= '0';
            internal_next_sm_mac_operation_mode <= "10";
            internal_next_mac_enable_reg_s_mask <= '0';
            internal_next_mac_subtraction_reg_a_b <= '0';
            internal_next_mac_sel_multiply_two_a_b <= '0';
            internal_next_mac_sel_reg_y_output <= '0';
            internal_next_sm_mac_write_enable_output <= '1';
            internal_next_mac_memory_double_mode <= '0';
            internal_next_mac_memory_only_write_mode <= '0';
            internal_next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_0 =>
            -- -- In case of size 1
            -- reg_a = a0_X; reg_b = a0_X; reg_acc = 0; Enable sign a,b; operation : a*b + acc;
            internal_next_sel_output_rom <= '1';
            internal_next_update_rom_address <= '1';
            internal_next_sel_load_new_rom_address <= '0';
            internal_next_sm_free_flag <= '0';
            internal_next_sm_rotation_size <= "11";
            internal_next_sm_circular_shift_enable <= '1';
            internal_next_sel_address_a <= '0';
            internal_next_sel_address_b_prime <= "00";
            internal_next_sm_specific_mac_address_a <= "000";
            internal_next_sm_specific_mac_address_b <= "000";
            internal_next_sm_specific_mac_address_o <= "000";
            internal_next_sm_specific_mac_next_address_o <= "001";
            internal_next_mac_enable_signed_a <= '1';
            internal_next_mac_enable_signed_b <= '1';
            internal_next_mac_sel_load_reg_a <= "00";
            internal_next_mac_clear_reg_b <= '0';
            internal_next_mac_clear_reg_acc <= '1';
            internal_next_mac_sel_shift_reg_o <= '0';
            internal_next_mac_enable_update_reg_s <= '0';
            internal_next_mac_sel_reg_s_reg_o_sign <= '0';
            internal_next_mac_reg_s_reg_o_positive <= '0';
            internal_next_sm_sign_a_mode <= '0';
            internal_next_sm_mac_operation_mode <= "10";
            internal_next_mac_enable_reg_s_mask <= '0';
            internal_next_mac_subtraction_reg_a_b <= '0';
            internal_next_mac_sel_multiply_two_a_b <= '0';
            internal_next_mac_sel_reg_y_output <= '0';
            internal_next_sm_mac_write_enable_output <= '0';
            internal_next_mac_memory_double_mode <= '0';
            internal_next_mac_memory_only_write_mode <= '0';
            internal_next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_5 =>
            -- -- In case of 2, 3, 4, 5, 6, 7, 8
            -- reg_a = a0_X; reg_b = a0_X; reg_acc = 0; operation : a*b + acc;
            internal_next_sel_output_rom <= '1';
            internal_next_update_rom_address <= '1';
            internal_next_sel_load_new_rom_address <= '0';
            internal_next_sm_free_flag <= '0';
            internal_next_sm_rotation_size <= "11";
            internal_next_sm_circular_shift_enable <= '1';
            internal_next_sel_address_a <= '0';
            internal_next_sel_address_b_prime <= "00";
            internal_next_sm_specific_mac_address_a <= "000";
            internal_next_sm_specific_mac_address_b <= "000";
            internal_next_sm_specific_mac_address_o <= "000";
            internal_next_sm_specific_mac_next_address_o <= "001";
            internal_next_mac_enable_signed_a <= '0';
            internal_next_mac_enable_signed_b <= '0';
            internal_next_mac_sel_load_reg_a <= "00";
            internal_next_mac_clear_reg_b <= '0';
            internal_next_mac_clear_reg_acc <= '1';
            internal_next_mac_sel_shift_reg_o <= '0';
            internal_next_mac_enable_update_reg_s <= '0';
            internal_next_mac_sel_reg_s_reg_o_sign <= '0';
            internal_next_mac_reg_s_reg_o_positive <= '0';
            internal_next_sm_sign_a_mode <= '0';
            internal_next_sm_mac_operation_mode <= "10";
            internal_next_mac_enable_reg_s_mask <= '0';
            internal_next_mac_subtraction_reg_a_b <= '0';
            internal_next_mac_sel_multiply_two_a_b <= '0';
            internal_next_mac_sel_reg_y_output <= '0';
            internal_next_sm_mac_write_enable_output <= '0';
            internal_next_mac_memory_double_mode <= '0';
            internal_next_mac_memory_only_write_mode <= '0';
            internal_next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_direct_0 =>
            -- -- In case of size 1
            -- reg_a = a0_X; reg_b = b0_X; reg_acc = 0; o0_0 = reg_o; Enable sign a,b; operation : b +/- a + acc;
            internal_next_sel_output_rom <= '1';
            internal_next_update_rom_address <= '1';
            internal_next_sel_load_new_rom_address <= '0';
            internal_next_sm_free_flag <= '0';
            internal_next_sm_rotation_size <= "10";
            internal_next_sm_circular_shift_enable <= '1';
            internal_next_sel_address_a <= '0';
            internal_next_sel_address_b_prime <= "00";
            internal_next_sm_specific_mac_address_a <= "000";
            internal_next_sm_specific_mac_address_b <= "000";
            internal_next_sm_specific_mac_address_o <= "000";
            internal_next_sm_specific_mac_next_address_o <= "001";
            internal_next_mac_enable_signed_a <= '1';
            internal_next_mac_enable_signed_b <= '1';
            internal_next_mac_sel_load_reg_a <= "00";
            internal_next_mac_clear_reg_b <= '0';
            internal_next_mac_clear_reg_acc <= '1';
            internal_next_mac_sel_shift_reg_o <= '0';
            internal_next_mac_enable_update_reg_s <= '0';
            internal_next_mac_sel_reg_s_reg_o_sign <= '0';
            internal_next_mac_reg_s_reg_o_positive <= '0';
            internal_next_sm_sign_a_mode <= '1';
            internal_next_sm_mac_operation_mode <= "00";
            internal_next_mac_enable_reg_s_mask <= '0';
            internal_next_mac_subtraction_reg_a_b <= '0';
            internal_next_mac_sel_multiply_two_a_b <= '0';
            internal_next_mac_sel_reg_y_output <= '0';
            internal_next_sm_mac_write_enable_output <= '1';
            internal_next_mac_memory_double_mode <= '0';
            internal_next_mac_memory_only_write_mode <= '0';
            internal_next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_direct_2 =>
            -- -- In case of size 2, 3, 4, 5, 6, 7, 8
            -- reg_a = a0_X; reg_b = b0_X; reg_acc = 0; o0_X = reg_o; operation : b +/- a + acc;
            internal_next_sel_output_rom <= '1';
            internal_next_update_rom_address <= '1';
            internal_next_sel_load_new_rom_address <= '0';
            internal_next_sm_free_flag <= '0';
            internal_next_sm_rotation_size <= "10";
            internal_next_sm_circular_shift_enable <= '1';
            internal_next_sel_address_a <= '0';
            internal_next_sel_address_b_prime <= "00";
            internal_next_sm_specific_mac_address_a <= "000";
            internal_next_sm_specific_mac_address_b <= "000";
            internal_next_sm_specific_mac_address_o <= "000";
            internal_next_sm_specific_mac_next_address_o <= "001";
            internal_next_mac_enable_signed_a <= '0';
            internal_next_mac_enable_signed_b <= '0';
            internal_next_mac_sel_load_reg_a <= "00";
            internal_next_mac_clear_reg_b <= '0';
            internal_next_mac_clear_reg_acc <= '1';
            internal_next_mac_sel_shift_reg_o <= '0';
            internal_next_mac_enable_update_reg_s <= '0';
            internal_next_mac_sel_reg_s_reg_o_sign <= '0';
            internal_next_mac_reg_s_reg_o_positive <= '0';
            internal_next_sm_sign_a_mode <= '1';
            internal_next_sm_mac_operation_mode <= "00";
            internal_next_mac_enable_reg_s_mask <= '0';
            internal_next_mac_subtraction_reg_a_b <= '0';
            internal_next_mac_sel_multiply_two_a_b <= '0';
            internal_next_mac_sel_reg_y_output <= '0';
            internal_next_sm_mac_write_enable_output <= '1';
            internal_next_mac_memory_double_mode <= '0';
            internal_next_mac_memory_only_write_mode <= '0';
            internal_next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_0 =>
            -- -- In case of size 1
            -- reg_a = a0_X; reg_b = 0; reg_acc = 0; Enable sign a,b; operation : b + a + acc;
            internal_next_sel_output_rom <= '1';
            internal_next_update_rom_address <= '1';
            internal_next_sel_load_new_rom_address <= '0';
            internal_next_sm_free_flag <= '0';
            internal_next_sm_rotation_size <= "10";
            internal_next_sm_circular_shift_enable <= '1';
            internal_next_sel_address_a <= '0';
            internal_next_sel_address_b_prime <= "10";
            internal_next_sm_specific_mac_address_a <= "000";
            internal_next_sm_specific_mac_address_b <= "000";
            internal_next_sm_specific_mac_address_o <= "000";
            internal_next_sm_specific_mac_next_address_o <= "001";
            internal_next_mac_enable_signed_a <= '1';
            internal_next_mac_enable_signed_b <= '1';
            internal_next_mac_sel_load_reg_a <= "00";
            internal_next_mac_clear_reg_b <= '1';
            internal_next_mac_clear_reg_acc <= '1';
            internal_next_mac_sel_shift_reg_o <= '0';
            internal_next_mac_enable_update_reg_s <= '0';
            internal_next_mac_sel_reg_s_reg_o_sign <= '0';
            internal_next_mac_reg_s_reg_o_positive <= '0';
            internal_next_sm_sign_a_mode <= '0';
            internal_next_sm_mac_operation_mode <= "01";
            internal_next_mac_enable_reg_s_mask <= '0';
            internal_next_mac_subtraction_reg_a_b <= '0';
            internal_next_mac_sel_multiply_two_a_b <= '0';
            internal_next_mac_sel_reg_y_output <= '0';
            internal_next_sm_mac_write_enable_output <= '0';
            internal_next_mac_memory_double_mode <= '0';
            internal_next_mac_memory_only_write_mode <= '0';
            internal_next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_5 =>
            -- -- In case of size 2
            -- reg_a = a1_X; reg_b = 0; reg_acc = 0; Enable sign a,b; operation : b + a + acc;
            internal_next_sel_output_rom <= '1';
            internal_next_update_rom_address <= '1';
            internal_next_sel_load_new_rom_address <= '0';
            internal_next_sm_free_flag <= '0';
            internal_next_sm_rotation_size <= "10";
            internal_next_sm_circular_shift_enable <= '1';
            internal_next_sel_address_a <= '0';
            internal_next_sel_address_b_prime <= "10";
            internal_next_sm_specific_mac_address_a <= "001";
            internal_next_sm_specific_mac_address_b <= "000";
            internal_next_sm_specific_mac_address_o <= "000";
            internal_next_sm_specific_mac_next_address_o <= "001";
            internal_next_mac_enable_signed_a <= '1';
            internal_next_mac_enable_signed_b <= '1';
            internal_next_mac_sel_load_reg_a <= "00";
            internal_next_mac_clear_reg_b <= '1';
            internal_next_mac_clear_reg_acc <= '1';
            internal_next_mac_sel_shift_reg_o <= '0';
            internal_next_mac_enable_update_reg_s <= '0';
            internal_next_mac_sel_reg_s_reg_o_sign <= '0';
            internal_next_mac_reg_s_reg_o_positive <= '0';
            internal_next_sm_sign_a_mode <= '0';
            internal_next_sm_mac_operation_mode <= "01";
            internal_next_mac_enable_reg_s_mask <= '0';
            internal_next_mac_subtraction_reg_a_b <= '0';
            internal_next_mac_sel_multiply_two_a_b <= '0';
            internal_next_mac_sel_reg_y_output <= '0';
            internal_next_sm_mac_write_enable_output <= '0';
            internal_next_mac_memory_double_mode <= '0';
            internal_next_mac_memory_only_write_mode <= '0';
            internal_next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_13 =>
            -- -- In case of size 3
            -- reg_a = a2_X; reg_b = 0; reg_acc = 0; Enable sign a,b; operation : b + a + acc;
            internal_next_sel_output_rom <= '1';
            internal_next_update_rom_address <= '1';
            internal_next_sel_load_new_rom_address <= '0';
            internal_next_sm_free_flag <= '0';
            internal_next_sm_rotation_size <= "10";
            internal_next_sm_circular_shift_enable <= '1';
            internal_next_sel_address_a <= '0';
            internal_next_sel_address_b_prime <= "10";
            internal_next_sm_specific_mac_address_a <= "010";
            internal_next_sm_specific_mac_address_b <= "010";
            internal_next_sm_specific_mac_address_o <= "010";
            internal_next_sm_specific_mac_next_address_o <= "011";
            internal_next_mac_enable_signed_a <= '1';
            internal_next_mac_enable_signed_b <= '1';
            internal_next_mac_sel_load_reg_a <= "00";
            internal_next_mac_clear_reg_b <= '1';
            internal_next_mac_clear_reg_acc <= '1';
            internal_next_mac_sel_shift_reg_o <= '0';
            internal_next_mac_enable_update_reg_s <= '0';
            internal_next_mac_sel_reg_s_reg_o_sign <= '0';
            internal_next_mac_reg_s_reg_o_positive <= '0';
            internal_next_sm_sign_a_mode <= '0';
            internal_next_sm_mac_operation_mode <= "01";
            internal_next_mac_enable_reg_s_mask <= '0';
            internal_next_mac_subtraction_reg_a_b <= '0';
            internal_next_mac_sel_multiply_two_a_b <= '0';
            internal_next_mac_sel_reg_y_output <= '0';
            internal_next_sm_mac_write_enable_output <= '0';
            internal_next_mac_memory_double_mode <= '0';
            internal_next_mac_memory_only_write_mode <= '0';
            internal_next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_24 =>
            -- -- In case of size 4
            -- reg_a = a3_X; reg_b = 0; reg_acc = 0; Enable sign a,b; operation : b + a + acc;
            internal_next_sel_output_rom <= '1';
            internal_next_update_rom_address <= '1';
            internal_next_sel_load_new_rom_address <= '0';
            internal_next_sm_free_flag <= '0';
            internal_next_sm_rotation_size <= "10";
            internal_next_sm_circular_shift_enable <= '1';
            internal_next_sel_address_a <= '0';
            internal_next_sel_address_b_prime <= "10";
            internal_next_sm_specific_mac_address_a <= "011";
            internal_next_sm_specific_mac_address_b <= "011";
            internal_next_sm_specific_mac_address_o <= "011";
            internal_next_sm_specific_mac_next_address_o <= "000";
            internal_next_mac_enable_signed_a <= '1';
            internal_next_mac_enable_signed_b <= '1';
            internal_next_mac_sel_load_reg_a <= "00";
            internal_next_mac_clear_reg_b <= '1';
            internal_next_mac_clear_reg_acc <= '1';
            internal_next_mac_sel_shift_reg_o <= '0';
            internal_next_mac_enable_update_reg_s <= '0';
            internal_next_mac_sel_reg_s_reg_o_sign <= '0';
            internal_next_mac_reg_s_reg_o_positive <= '0';
            internal_next_sm_sign_a_mode <= '0';
            internal_next_sm_mac_operation_mode <= "01";
            internal_next_mac_enable_reg_s_mask <= '0';
            internal_next_mac_subtraction_reg_a_b <= '0';
            internal_next_mac_sel_multiply_two_a_b <= '0';
            internal_next_mac_sel_reg_y_output <= '0';
            internal_next_sm_mac_write_enable_output <= '0';
            internal_next_mac_memory_double_mode <= '0';
            internal_next_mac_memory_only_write_mode <= '0';
            internal_next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_38 =>
            -- -- In case of size 5
            -- reg_a = a4_X; reg_b = 0; reg_acc = 0; Enable sign a,b; operation : b + a + acc;
            internal_next_sel_output_rom <= '1';
            internal_next_update_rom_address <= '1';
            internal_next_sel_load_new_rom_address <= '0';
            internal_next_sm_free_flag <= '0';
            internal_next_sm_rotation_size <= "10";
            internal_next_sm_circular_shift_enable <= '1';
            internal_next_sel_address_a <= '0';
            internal_next_sel_address_b_prime <= "10";
            internal_next_sm_specific_mac_address_a <= "100";
            internal_next_sm_specific_mac_address_b <= "100";
            internal_next_sm_specific_mac_address_o <= "100";
            internal_next_sm_specific_mac_next_address_o <= "101";
            internal_next_mac_enable_signed_a <= '1';
            internal_next_mac_enable_signed_b <= '1';
            internal_next_mac_sel_load_reg_a <= "00";
            internal_next_mac_clear_reg_b <= '1';
            internal_next_mac_clear_reg_acc <= '1';
            internal_next_mac_sel_shift_reg_o <= '0';
            internal_next_mac_enable_update_reg_s <= '0';
            internal_next_mac_sel_reg_s_reg_o_sign <= '0';
            internal_next_mac_reg_s_reg_o_positive <= '0';
            internal_next_sm_sign_a_mode <= '0';
            internal_next_sm_mac_operation_mode <= "01";
            internal_next_mac_enable_reg_s_mask <= '0';
            internal_next_mac_subtraction_reg_a_b <= '0';
            internal_next_mac_sel_multiply_two_a_b <= '0';
            internal_next_mac_sel_reg_y_output <= '0';
            internal_next_sm_mac_write_enable_output <= '0';
            internal_next_mac_memory_double_mode <= '0';
            internal_next_mac_memory_only_write_mode <= '0';
            internal_next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_55 =>
            -- -- In case of size 6
            -- reg_a = a5_X; reg_b = 0; reg_acc = 0; Enable sign a,b; operation : b + a + acc;
            internal_next_sel_output_rom <= '1';
            internal_next_update_rom_address <= '1';
            internal_next_sel_load_new_rom_address <= '0';
            internal_next_sm_free_flag <= '0';
            internal_next_sm_rotation_size <= "10";
            internal_next_sm_circular_shift_enable <= '1';
            internal_next_sel_address_a <= '0';
            internal_next_sel_address_b_prime <= "10";
            internal_next_sm_specific_mac_address_a <= "101";
            internal_next_sm_specific_mac_address_b <= "101";
            internal_next_sm_specific_mac_address_o <= "101";
            internal_next_sm_specific_mac_next_address_o <= "110";
            internal_next_mac_enable_signed_a <= '1';
            internal_next_mac_enable_signed_b <= '1';
            internal_next_mac_sel_load_reg_a <= "00";
            internal_next_mac_clear_reg_b <= '1';
            internal_next_mac_clear_reg_acc <= '1';
            internal_next_mac_sel_shift_reg_o <= '0';
            internal_next_mac_enable_update_reg_s <= '0';
            internal_next_mac_sel_reg_s_reg_o_sign <= '0';
            internal_next_mac_reg_s_reg_o_positive <= '0';
            internal_next_sm_sign_a_mode <= '0';
            internal_next_sm_mac_operation_mode <= "01";
            internal_next_mac_enable_reg_s_mask <= '0';
            internal_next_mac_subtraction_reg_a_b <= '0';
            internal_next_mac_sel_multiply_two_a_b <= '0';
            internal_next_mac_sel_reg_y_output <= '0';
            internal_next_sm_mac_write_enable_output <= '0';
            internal_next_mac_memory_double_mode <= '0';
            internal_next_mac_memory_only_write_mode <= '0';
            internal_next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_75 =>
            -- -- In case of size 7
            -- reg_a = a6_X; reg_b = 0; reg_acc = 0; Enable sign a,b; operation : b + a + acc;
            internal_next_sel_output_rom <= '1';
            internal_next_update_rom_address <= '1';
            internal_next_sel_load_new_rom_address <= '0';
            internal_next_sm_free_flag <= '0';
            internal_next_sm_rotation_size <= "10";
            internal_next_sm_circular_shift_enable <= '1';
            internal_next_sel_address_a <= '0';
            internal_next_sel_address_b_prime <= "10";
            internal_next_sm_specific_mac_address_a <= "110";
            internal_next_sm_specific_mac_address_b <= "110";
            internal_next_sm_specific_mac_address_o <= "110";
            internal_next_sm_specific_mac_next_address_o <= "111";
            internal_next_mac_enable_signed_a <= '1';
            internal_next_mac_enable_signed_b <= '1';
            internal_next_mac_sel_load_reg_a <= "00";
            internal_next_mac_clear_reg_b <= '1';
            internal_next_mac_clear_reg_acc <= '1';
            internal_next_mac_sel_shift_reg_o <= '0';
            internal_next_mac_enable_update_reg_s <= '0';
            internal_next_mac_sel_reg_s_reg_o_sign <= '0';
            internal_next_mac_reg_s_reg_o_positive <= '0';
            internal_next_sm_sign_a_mode <= '0';
            internal_next_sm_mac_operation_mode <= "01";
            internal_next_mac_enable_reg_s_mask <= '0';
            internal_next_mac_subtraction_reg_a_b <= '0';
            internal_next_mac_sel_multiply_two_a_b <= '0';
            internal_next_mac_sel_reg_y_output <= '0';
            internal_next_sm_mac_write_enable_output <= '0';
            internal_next_mac_memory_double_mode <= '0';
            internal_next_mac_memory_only_write_mode <= '0';
            internal_next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_98 =>
            -- -- In case of size 8
            -- reg_a = a7_X; reg_b = 0; reg_acc = 0; Enable sign a,b; operation : b + a + acc;
            internal_next_sel_output_rom <= '1';
            internal_next_update_rom_address <= '1';
            internal_next_sel_load_new_rom_address <= '0';
            internal_next_sm_free_flag <= '0';
            internal_next_sm_rotation_size <= "10";
            internal_next_sm_circular_shift_enable <= '1';
            internal_next_sel_address_a <= '0';
            internal_next_sel_address_b_prime <= "10";
            internal_next_sm_specific_mac_address_a <= "111";
            internal_next_sm_specific_mac_address_b <= "111";
            internal_next_sm_specific_mac_address_o <= "111";
            internal_next_sm_specific_mac_next_address_o <= "000";
            internal_next_mac_enable_signed_a <= '1';
            internal_next_mac_enable_signed_b <= '1';
            internal_next_mac_sel_load_reg_a <= "00";
            internal_next_mac_clear_reg_b <= '1';
            internal_next_mac_clear_reg_acc <= '1';
            internal_next_mac_sel_shift_reg_o <= '0';
            internal_next_mac_enable_update_reg_s <= '0';
            internal_next_mac_sel_reg_s_reg_o_sign <= '0';
            internal_next_mac_reg_s_reg_o_positive <= '0';
            internal_next_sm_sign_a_mode <= '0';
            internal_next_sm_mac_operation_mode <= "01";
            internal_next_mac_enable_reg_s_mask <= '0';
            internal_next_mac_subtraction_reg_a_b <= '0';
            internal_next_mac_sel_multiply_two_a_b <= '0';
            internal_next_mac_sel_reg_y_output <= '0';
            internal_next_sm_mac_write_enable_output <= '0';
            internal_next_mac_memory_double_mode <= '0';
            internal_next_mac_memory_only_write_mode <= '0';
            internal_next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_0 =>
            -- Operands size 1
            -- reg_a = a0_X; reg_b = b0_X; reg_acc = 0; o0_X = reg_o; Enable sign a,b; operation : b +/- a + acc;
            internal_next_sel_output_rom <= '1';
            internal_next_update_rom_address <= '1';
            internal_next_sel_load_new_rom_address <= '0';
            internal_next_sm_free_flag <= '0';
            internal_next_sm_rotation_size <= "10";
            internal_next_sm_circular_shift_enable <= '1';
            internal_next_sel_address_a <= '0';
            internal_next_sel_address_b_prime <= "00";
            internal_next_sm_specific_mac_address_a <= "000";
            internal_next_sm_specific_mac_address_b <= "000";
            internal_next_sm_specific_mac_address_o <= "000";
            internal_next_sm_specific_mac_next_address_o <= "001";
            internal_next_mac_enable_signed_a <= '1';
            internal_next_mac_enable_signed_b <= '1';
            internal_next_mac_sel_load_reg_a <= "00";
            internal_next_mac_clear_reg_b <= '0';
            internal_next_mac_clear_reg_acc <= '1';
            internal_next_mac_sel_shift_reg_o <= '0';
            internal_next_mac_enable_update_reg_s <= '0';
            internal_next_mac_sel_reg_s_reg_o_sign <= '0';
            internal_next_mac_reg_s_reg_o_positive <= '0';
            internal_next_sm_sign_a_mode <= '1';
            internal_next_sm_mac_operation_mode <= "01";
            internal_next_mac_enable_reg_s_mask <= '0';
            internal_next_mac_subtraction_reg_a_b <= '0';
            internal_next_mac_sel_multiply_two_a_b <= '0';
            internal_next_mac_sel_reg_y_output <= '0';
            internal_next_sm_mac_write_enable_output <= '1';
            internal_next_mac_memory_double_mode <= '0';
            internal_next_mac_memory_only_write_mode <= '0';
            internal_next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_with_reduction_5 =>
            -- -- In case of sizes 2, 3, 4, 5, 6, 7, 8
            -- reg_a = a0_X; reg_b = b0_X; reg_acc = 0; o0_X = reg_o; operation : b +/- a + acc;
            internal_next_sel_output_rom <= '1';
            internal_next_update_rom_address <= '1';
            internal_next_sel_load_new_rom_address <= '0';
            internal_next_sm_free_flag <= '0';
            internal_next_sm_rotation_size <= "10";
            internal_next_sm_circular_shift_enable <= '1';
            internal_next_sel_address_a <= '0';
            internal_next_sel_address_b_prime <= "00";
            internal_next_sm_specific_mac_address_a <= "000";
            internal_next_sm_specific_mac_address_b <= "000";
            internal_next_sm_specific_mac_address_o <= "000";
            internal_next_sm_specific_mac_next_address_o <= "001";
            internal_next_mac_enable_signed_a <= '0';
            internal_next_mac_enable_signed_b <= '0';
            internal_next_mac_sel_load_reg_a <= "00";
            internal_next_mac_clear_reg_b <= '0';
            internal_next_mac_clear_reg_acc <= '1';
            internal_next_mac_sel_shift_reg_o <= '0';
            internal_next_mac_enable_update_reg_s <= '0';
            internal_next_mac_sel_reg_s_reg_o_sign <= '0';
            internal_next_mac_reg_s_reg_o_positive <= '0';
            internal_next_sm_sign_a_mode <= '1';
            internal_next_sm_mac_operation_mode <= "00";
            internal_next_mac_enable_reg_s_mask <= '0';
            internal_next_mac_subtraction_reg_a_b <= '0';
            internal_next_mac_sel_multiply_two_a_b <= '0';
            internal_next_mac_sel_reg_y_output <= '0';
            internal_next_sm_mac_write_enable_output <= '1';
            internal_next_mac_memory_double_mode <= '0';
            internal_next_mac_memory_only_write_mode <= '0';
            internal_next_base_address_generator_o_increment_previous_address <= '0';
        when instruction_execution =>
            internal_next_sel_output_rom <= '1';
            internal_next_update_rom_address <= '1';
            internal_next_sel_load_new_rom_address <= '0';
            internal_next_sm_free_flag <= '0';
            internal_next_sm_rotation_size <= "11";
            internal_next_sm_circular_shift_enable <= '1';
            internal_next_sel_address_a <= '0';
            internal_next_sel_address_b_prime <= "00";
            internal_next_sm_specific_mac_address_a <= "000";
            internal_next_sm_specific_mac_address_b <= "000";
            internal_next_sm_specific_mac_address_o <= "000";
            internal_next_sm_specific_mac_next_address_o <= "001";
            internal_next_mac_enable_signed_a <= '0';
            internal_next_mac_enable_signed_b <= '0';
            internal_next_mac_sel_load_reg_a <= "11";
            internal_next_mac_clear_reg_b <= '1';
            internal_next_mac_clear_reg_acc <= '1';
            internal_next_mac_sel_shift_reg_o <= '0';
            internal_next_mac_enable_update_reg_s <= '0';
            internal_next_mac_sel_reg_s_reg_o_sign <= '0';
            internal_next_mac_reg_s_reg_o_positive <= '0';
            internal_next_sm_sign_a_mode <= '0';
            internal_next_sm_mac_operation_mode <= "10";
            internal_next_mac_enable_reg_s_mask <= '0';
            internal_next_mac_subtraction_reg_a_b <= '0';
            internal_next_mac_sel_multiply_two_a_b <= '0';
            internal_next_mac_sel_reg_y_output <= '0';
            internal_next_sm_mac_write_enable_output <= '0';
            internal_next_mac_memory_double_mode <= '0';
            internal_next_mac_memory_only_write_mode <= '0';
            internal_next_base_address_generator_o_increment_previous_address <= '0';
    end case;
end process;

update_state : process(actual_state, instruction_type, operands_size, instruction_values_valid, prime_line_equal_one, ultimate_instruction, reg_rom_last_state)
begin
case (actual_state) is
        when reset =>
            next_state <= decode_instruction;
        when decode_instruction =>
            next_state <= decode_instruction;
            if(instruction_values_valid = '1') then
                if(instruction_type = "0000") then
                    if(operands_size = "000") then
                        next_state <= multiplication_direct_0;
                    else
                        next_state <= multiplication_direct_2;
                    end if;
                elsif(instruction_type = "0001") then
                    if(operands_size = "000") then
                        next_state <= square_direct_0;
                    else
                        next_state <= square_direct_2;
                    end if;
                elsif(instruction_type = "0010") then
                    case (prime_line_equal_one) is
                        when "00" =>
                            if(operands_size = "000") then
                                next_state <= multiplication_with_reduction_0;
                            else
                                next_state <= multiplication_with_reduction_5;
                            end if;
                        when "01" =>
                            if(operands_size = "000") then
                                next_state <= multiplication_with_reduction_special_prime_1_0;
                            else
                                next_state <= multiplication_with_reduction_special_prime_1_3;
                            end if;
                        when "10" =>
                            next_state <= multiplication_with_reduction_special_prime_2_0;
                        when "11" =>
                            next_state <= multiplication_with_reduction_special_prime_3_0;
                        when others =>
                            next_state <= decode_instruction;
                    end case;
                elsif(instruction_type = "0011") then
                    case (prime_line_equal_one) is
                        when "00" =>
                            if(operands_size = "000") then
                                next_state <= square_with_reduction_0;
                            else
                                next_state <= square_with_reduction_5;
                            end if;
                        when "01" =>
                            if(operands_size = "000") then
                                next_state <= square_with_reduction_special_prime_1_0;
                            else
                                next_state <= square_with_reduction_special_prime_1_3;
                            end if;
                        when "10" =>
                            next_state <= square_with_reduction_special_prime_2_0;
                        when "11" =>
                            next_state <= square_with_reduction_special_prime_3_0;
                        when others =>
                            next_state <= decode_instruction;
                    end case;
                elsif(instruction_type = "0100") then
                    if(operands_size = "000") then
                        next_state <= addition_subtraction_direct_0;
                    else
                        next_state <= addition_subtraction_direct_2;
                    end if;
                elsif(instruction_type = "0101") then
                    if(operands_size = "000") then
                        next_state <= iterative_modular_reduction_0;
                    elsif(operands_size = "001") then
                        next_state <= iterative_modular_reduction_5;
                    elsif(operands_size = "010") then
                        next_state <= iterative_modular_reduction_13;
                    elsif(operands_size = "011") then
                        next_state <= iterative_modular_reduction_24;
                    elsif(operands_size = "100") then
                        next_state <= iterative_modular_reduction_38;
                    elsif(operands_size = "101") then
                        next_state <= iterative_modular_reduction_55;
                    elsif(operands_size = "110") then
                        next_state <= iterative_modular_reduction_75;
                    else
                        next_state <= iterative_modular_reduction_98;
                    end if;
                elsif(instruction_type = "0110") then
                    if(operands_size = "000") then
                        next_state <= addition_subtraction_with_reduction_0;
                    else
                        next_state <= addition_subtraction_with_reduction_5;
                    end if;
                end if;
            end if;
        when multiplication_direct_0 =>
            next_state <= multiplication_direct_0;
            if(ultimate_instruction = '1') then
                next_state <= instruction_execution;
            end if;
        when multiplication_direct_2 =>
            next_state <= multiplication_direct_2;
            if(ultimate_instruction = '1') then
                next_state <= instruction_execution;
            end if;
        when square_direct_0 =>
            next_state <= square_direct_0;
            if(ultimate_instruction = '1') then
                next_state <= instruction_execution;
            end if;
        when square_direct_2 =>
            next_state <= square_direct_2;
            if(ultimate_instruction = '1') then
                next_state <= instruction_execution;
            end if;
        when multiplication_with_reduction_special_prime_1_0 =>
            next_state <= multiplication_with_reduction_special_prime_1_0;
            if(ultimate_instruction = '1') then
                next_state <= instruction_execution;
            end if;
        when multiplication_with_reduction_special_prime_1_3 =>
            next_state <= multiplication_with_reduction_special_prime_1_3;
            if(ultimate_instruction = '1') then
                next_state <= instruction_execution;
            end if;
        when multiplication_with_reduction_special_prime_2_0 =>
            next_state <= multiplication_with_reduction_special_prime_2_0;
            if(ultimate_instruction = '1') then
                next_state <= instruction_execution;
            end if;
        when multiplication_with_reduction_special_prime_3_0 =>
            next_state <= multiplication_with_reduction_special_prime_3_0;
            if(ultimate_instruction = '1') then
                next_state <= instruction_execution;
            end if;
        when multiplication_with_reduction_0 =>
            next_state <= multiplication_with_reduction_0;
            if(ultimate_instruction = '1') then
                next_state <= instruction_execution;
            end if;
        when multiplication_with_reduction_5 =>
            next_state <= multiplication_with_reduction_5;
            if(ultimate_instruction = '1') then
                next_state <= instruction_execution;
            end if;
        when square_with_reduction_special_prime_1_0 =>
            next_state <= square_with_reduction_special_prime_1_0;
            if(ultimate_instruction = '1') then
                next_state <= instruction_execution;
            end if;
        when square_with_reduction_special_prime_1_3 =>
            next_state <= square_with_reduction_special_prime_1_3;
            if(ultimate_instruction = '1') then
                next_state <= instruction_execution;
            end if;
        when square_with_reduction_special_prime_2_0 =>
            next_state <= square_with_reduction_special_prime_2_0;
            if(ultimate_instruction = '1') then
                next_state <= instruction_execution;
            end if;
        when square_with_reduction_special_prime_3_0 =>
            next_state <= square_with_reduction_special_prime_3_0;
            if(ultimate_instruction = '1') then
                next_state <= instruction_execution;
            end if;
        when square_with_reduction_0 =>
            next_state <= square_with_reduction_0;
            if(ultimate_instruction = '1') then
                next_state <= instruction_execution;
            end if;
        when square_with_reduction_5 =>
            next_state <= square_with_reduction_5;
            if(ultimate_instruction = '1') then
                next_state <= instruction_execution;
            end if;
        when addition_subtraction_direct_0 =>
            next_state <= addition_subtraction_direct_0;
            if(ultimate_instruction = '1') then
                next_state <= instruction_execution;
            end if;
        when addition_subtraction_direct_2 =>
            next_state <= addition_subtraction_direct_2;
            if(ultimate_instruction = '1') then
                next_state <= instruction_execution;
            end if;
        when iterative_modular_reduction_0 =>
            next_state <= iterative_modular_reduction_0;
            if(ultimate_instruction = '1') then
                next_state <= instruction_execution;
            end if;
        when iterative_modular_reduction_5 =>
            next_state <= iterative_modular_reduction_5;
            if(ultimate_instruction = '1') then
                next_state <= instruction_execution;
            end if;
        when iterative_modular_reduction_13 =>
            next_state <= iterative_modular_reduction_13;
            if(ultimate_instruction = '1') then
                next_state <= instruction_execution;
            end if;
        when iterative_modular_reduction_24 =>
            next_state <= iterative_modular_reduction_24;
            if(ultimate_instruction = '1') then
                next_state <= instruction_execution;
            end if;
        when iterative_modular_reduction_38 =>
            next_state <= iterative_modular_reduction_38;
            if(ultimate_instruction = '1') then
                next_state <= instruction_execution;
            end if;
        when iterative_modular_reduction_55 =>
            next_state <= iterative_modular_reduction_55;
            if(ultimate_instruction = '1') then
                next_state <= instruction_execution;
            end if;
        when iterative_modular_reduction_75 =>
            next_state <= iterative_modular_reduction_75;
            if(ultimate_instruction = '1') then
                next_state <= instruction_execution;
            end if;
        when iterative_modular_reduction_98 =>
            next_state <= iterative_modular_reduction_98;
            if(ultimate_instruction = '1') then
                next_state <= instruction_execution;
            end if;
        when addition_subtraction_with_reduction_0 =>
            next_state <= addition_subtraction_with_reduction_0;
            if(ultimate_instruction = '1') then
                next_state <= instruction_execution;
            end if;
        when addition_subtraction_with_reduction_5 =>
            next_state <= addition_subtraction_with_reduction_5;
            if(ultimate_instruction = '1') then
                next_state <= instruction_execution;
            end if;
        when instruction_execution =>
            next_state <= instruction_execution;
            if((ultimate_instruction = '1') and (reg_rom_last_state = '1')) then
                next_state <= decode_instruction;
            end if;
end case;
end process;

process(clk)
begin
    if(rising_edge(clk)) then
        if(rstn = '0') then
            ultimate_instruction <= '0';
        else
            ultimate_instruction <= penultimate_operation;
        end if;
    end if;
end process;

adder_a <= unsigned(rom_state_machine_address);
adder_b <= resize(unsigned(rom_next_operation_same_operand_size), adder_b'length) when (rom_current_operand_size = operands_size) else unsigned(rom_next_operation_different_operand_size);

adder_o <= adder_a + resize(adder_b, adder_o'length);

process(clk)
begin
    if (rising_edge(clk)) then
        rom_state_machine_address <= rom_state_machine_next_address;
    end if;
end process;

process(rom_state_machine_address, internal_update_rom_address, internal_sel_load_new_rom_address, instruction_values_valid, instruction_type, operands_size, prime_line_equal_one, penultimate_operation, adder_o)
begin
    if(internal_update_rom_address = '0') then
        rom_state_machine_next_address <= rom_state_machine_address;
    else
        if(internal_sel_load_new_rom_address = '1') then
            if(instruction_values_valid = '1') then
                if(instruction_type = "0000") then
                    if(operands_size = "000") then
                        rom_state_machine_next_address <= first_state_multiplication_direct_operand_size_1;
                    else
                        rom_state_machine_next_address <= first_state_multiplication_direct_operand_size_2_3_4_5_6_7_8;
                    end if;
                elsif(instruction_type = "0001") then
                    if(operands_size = "000") then
                        rom_state_machine_next_address <= first_state_square_direct_operand_size_1;
                    else
                        rom_state_machine_next_address <= first_state_square_direct_operand_size_2_3_4_5_6_7_8;
                    end if;
                elsif(instruction_type = "0010") then
                    case (prime_line_equal_one) is
                        when "00" =>
                            if(operands_size = "000") then
                                rom_state_machine_next_address <= first_state_multiplication_with_reduction_operand_size_1;
                            else
                                rom_state_machine_next_address <= first_state_multiplication_with_reduction_operand_size_2_3_4_5_6_7_8;
                            end if;
                        when "01" =>
                            if(operands_size = "000") then
                                rom_state_machine_next_address <= first_state_multiplication_with_reduction_special_prime_1_operand_size_1;
                            else
                                rom_state_machine_next_address <= first_state_multiplication_with_reduction_special_prime_1_operand_size_2_3_4_5_6_7_8;
                            end if;
                        when "10" =>
                            rom_state_machine_next_address <= first_state_multiplication_with_reduction_special_prime_2_operand_size_2_3_4_5_6_7_8;
                        when "11" =>
                            rom_state_machine_next_address <= first_state_multiplication_with_reduction_special_prime_3_operand_size_3_4_5_6_7_8;
                        when others =>
                            rom_state_machine_next_address <= rom_state_machine_address;
                    end case;
                elsif(instruction_type = "0011") then
                    case (prime_line_equal_one) is
                        when "00" =>
                            if(operands_size = "000") then
                                rom_state_machine_next_address <= first_state_square_with_reduction_operand_size_1;
                            else
                                rom_state_machine_next_address <= first_state_square_with_reduction_operand_size_2_3_4_5_6_7_8;
                            end if;
                        when "01" =>
                            if(operands_size = "000") then
                                rom_state_machine_next_address <= first_state_square_with_reduction_special_prime_1_operand_size_1;
                            else
                                rom_state_machine_next_address <= first_state_square_with_reduction_special_prime_1_operand_size_2_3_4_5_6_7_8;
                            end if;
                        when "10" =>
                            rom_state_machine_next_address <= first_state_square_with_reduction_special_prime_2_operand_size_2_3_4_5_6_7_8;
                        when "11" =>
                            rom_state_machine_next_address <= first_state_square_with_reduction_special_prime_3_operand_size_3_4_5_6_7_8;
                        when others =>
                            rom_state_machine_next_address <= rom_state_machine_address;
                    end case;
                elsif(instruction_type = "0100") then
                    if(operands_size = "000") then
                        rom_state_machine_next_address <= first_state_addition_subtraction_direct_operand_size_1;
                    else
                        rom_state_machine_next_address <= first_state_addition_subtraction_direct_operand_size_2_3_4_5_6_7_8;
                    end if;
                elsif(instruction_type = "0101") then
                    if(operands_size = "000") then
                        rom_state_machine_next_address <= first_state_iterative_modular_reduction_operand_size_1;
                    elsif(operands_size = "001") then
                        rom_state_machine_next_address <= first_state_iterative_modular_reduction_operand_size_2;
                    elsif(operands_size = "010") then
                        rom_state_machine_next_address <= first_state_iterative_modular_reduction_operand_size_3;
                    elsif(operands_size = "011") then
                        rom_state_machine_next_address <= first_state_iterative_modular_reduction_operand_size_4;
                    elsif(operands_size = "100") then
                        rom_state_machine_next_address <= first_state_iterative_modular_reduction_operand_size_5;
                    elsif(operands_size = "101") then
                        rom_state_machine_next_address <= first_state_iterative_modular_reduction_operand_size_6;
                    elsif(operands_size = "110") then
                        rom_state_machine_next_address <= first_state_iterative_modular_reduction_operand_size_7;
                    else
                        rom_state_machine_next_address <= first_state_iterative_modular_reduction_operand_size_8;
                    end if;
                elsif(instruction_type = "0110") then
                    if(operands_size = "000") then
                        rom_state_machine_next_address <= first_state_addition_subtraction_with_reduction_operand_size_1;
                    else
                        rom_state_machine_next_address <= first_state_addition_subtraction_with_reduction_operand_size_2_3_4_5_6_7_8;
                    end if;
                else
                    rom_state_machine_next_address <= rom_state_machine_address;
                end if;
            else
                rom_state_machine_next_address <= rom_state_machine_address;
            end if;
        elsif(penultimate_operation = '1') then
            rom_state_machine_next_address <= std_logic_vector(adder_o);
        else
            rom_state_machine_next_address <= rom_state_machine_address;
        end if;
    end if;
end process;

rom_state_machine_output <= rom_state_machine(to_integer(to_01(unsigned(rom_state_machine_address))));

rom_sm_rotation_size <= rom_state_machine_output(1 downto 0);
rom_sel_address_a <= rom_state_machine_output(2);
rom_sel_address_b_prime <= rom_state_machine_output(4 downto 3);
rom_sm_specific_mac_address_a <= rom_state_machine_output(7 downto 5);
rom_sm_specific_mac_address_b <= rom_state_machine_output(10 downto 8);
rom_sm_specific_mac_address_o <= rom_state_machine_output(13 downto 11);
rom_sm_specific_mac_next_address_o <= rom_state_machine_output(16 downto 14);
rom_mac_enable_signed_a <= rom_state_machine_output(17);
rom_mac_enable_signed_b <= rom_state_machine_output(18);
rom_mac_sel_load_reg_a <= rom_state_machine_output(20 downto 19);
rom_mac_clear_reg_b <= rom_state_machine_output(21);
rom_mac_clear_reg_acc <= rom_state_machine_output(22);
rom_mac_sel_shift_reg_o <= rom_state_machine_output(23);
rom_mac_enable_update_reg_s <= rom_state_machine_output(24);
rom_mac_sel_reg_s_reg_o_sign <= rom_state_machine_output(25);
rom_mac_reg_s_reg_o_positive <= rom_state_machine_output(26);
rom_sm_sign_a_mode <= rom_state_machine_output(27);
rom_sm_mac_operation_mode <= rom_state_machine_output(29 downto 28);
rom_mac_enable_reg_s_mask <= rom_state_machine_output(30);
rom_mac_subtraction_reg_a_b <= rom_state_machine_output(31);
rom_mac_sel_multiply_two_a_b <= rom_state_machine_output(32);
rom_mac_sel_reg_y_output <= rom_state_machine_output(33);
rom_sm_mac_write_enable_output <= rom_state_machine_output(34);
rom_mac_memory_double_mode <= rom_state_machine_output(35);
rom_mac_memory_only_write_mode <= rom_state_machine_output(36);
rom_base_address_generator_o_increment_previous_address <= rom_state_machine_output(37);

rom_last_state <= rom_state_machine_output(38);
rom_current_operand_size <= rom_state_machine_output(41 downto 39);
rom_next_operation_same_operand_size <= rom_state_machine_output(46 downto 42);
rom_next_operation_different_operand_size <= rom_state_machine_output(53 downto 47);

process(clk)
begin
    if(rising_edge(clk)) then
        if(rstn = '0') then
            reg_rom_last_state <= '0';
        else
            reg_rom_last_state <= rom_last_state;
        end if;
    end if;
end process;

sm_rotation_size <= internal_sm_rotation_size;
sm_circular_shift_enable <= internal_sm_circular_shift_enable;
sel_address_a <= internal_sel_address_a;
sel_address_b_prime <= internal_sel_address_b_prime;
sm_specific_mac_address_a <= internal_sm_specific_mac_address_a;
sm_specific_mac_address_b <= internal_sm_specific_mac_address_b;
sm_specific_mac_address_o <= internal_sm_specific_mac_address_o;
sm_specific_mac_next_address_o <= internal_sm_specific_mac_next_address_o;
mac_enable_signed_a <= internal_mac_enable_signed_a;
mac_enable_signed_b <= internal_mac_enable_signed_b;
mac_sel_load_reg_a <= internal_mac_sel_load_reg_a;
mac_clear_reg_b <= internal_mac_clear_reg_b;
mac_clear_reg_acc <= internal_mac_clear_reg_acc;
mac_sel_shift_reg_o <= internal_mac_sel_shift_reg_o;
mac_enable_update_reg_s <= internal_mac_enable_update_reg_s;
mac_sel_reg_s_reg_o_sign <= internal_mac_sel_reg_s_reg_o_sign;
mac_reg_s_reg_o_positive <= internal_mac_reg_s_reg_o_positive;
sm_sign_a_mode <= internal_sm_sign_a_mode;
sm_mac_operation_mode <= internal_sm_mac_operation_mode;
mac_enable_reg_s_mask <= internal_mac_enable_reg_s_mask;
mac_subtraction_reg_a_b <= internal_mac_subtraction_reg_a_b;
mac_sel_multiply_two_a_b <= internal_mac_sel_multiply_two_a_b;
mac_sel_reg_y_output <= internal_mac_sel_reg_y_output;
sm_mac_write_enable_output <= internal_sm_mac_write_enable_output;
mac_memory_double_mode <= internal_mac_memory_double_mode;
mac_memory_only_write_mode <= internal_mac_memory_only_write_mode;
base_address_generator_o_increment_previous_address <= internal_base_address_generator_o_increment_previous_address;
sm_free_flag <= internal_sm_free_flag;

end compact_memory_based_v3;