--
-- Implementation by Pedro Maat C. Massolino, hereby denoted as "the implementer".
--
-- To the extent possible under law, the implementer has waived all copyright
-- and related or neighboring rights to the source code in this file.
-- http://creativecommons.org/publicdomain/zero/1.0/
--
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity carmela_state_machine_v256 is
    Port (
        clk : in std_logic;
        rstn : in std_logic;
        instruction_values_valid : in std_logic;
        instruction_type : in std_logic_vector(3 downto 0);
        operands_size : in std_logic_vector(1 downto 0);
        prime_line_equal_one : in std_logic;
        penultimate_operation : in std_logic;
        sm_rotation_size : out std_logic_vector(1 downto 0);
        sm_circular_shift_enable : out std_logic;
        sel_address_a : out std_logic;
        sel_address_b_prime : out std_logic_vector(1 downto 0);
        sm_specific_mac_address_a : out std_logic_vector(1 downto 0);
        sm_specific_mac_address_b : out std_logic_vector(1 downto 0);
        sm_specific_mac_address_o : out std_logic_vector(1 downto 0);
        sm_specific_mac_next_address_o : out std_logic_vector(1 downto 0);
        mac_enable_signed_a : out std_logic;
        mac_enable_signed_b : out std_logic;
        mac_sel_load_reg_a : out std_logic_vector(1 downto 0);
        mac_clear_reg_b : out std_logic;
        mac_clear_reg_acc : out std_logic;
        mac_sel_shift_reg_o : out std_logic;
        mac_enable_update_reg_s : out std_logic;
        mac_sel_reg_s_reg_o_sign : out std_logic;
        mac_reg_s_reg_o_positive : out std_logic;
        sm_sign_a_mode : out std_logic;
        sm_mac_operation_mode : out std_logic_vector(1 downto 0);
        mac_enable_reg_s_mask : out std_logic;
        mac_subtraction_reg_a_b : out std_logic;
        mac_sel_multiply_two_a_b : out std_logic;
        mac_sel_reg_y_output : out std_logic;
        sm_mac_write_enable_output : out std_logic;
        mac_memory_double_mode : out std_logic;
        mac_memory_only_write_mode : out std_logic;
        base_address_generator_o_increment_previous_address : out std_logic;
        sm_free_flag : out std_logic
    );
end carmela_state_machine_v256;

architecture behavioral of carmela_state_machine_v256 is

type state is (reset, decode_instruction,
-- 0000 multiplication with no reduction
multiplication_direct_0, multiplication_direct_2, multiplication_direct_3, multiplication_direct_4, multiplication_direct_5, multiplication_direct_7, multiplication_direct_8, multiplication_direct_9, multiplication_direct_10, multiplication_direct_11, multiplication_direct_12, multiplication_direct_13, multiplication_direct_14, multiplication_direct_16, multiplication_direct_17, multiplication_direct_18, multiplication_direct_19, multiplication_direct_20, multiplication_direct_21, multiplication_direct_22, multiplication_direct_23, multiplication_direct_24, multiplication_direct_25, multiplication_direct_26, multiplication_direct_27,
-- 0001 square with no reduction
square_direct_0, square_direct_2, square_direct_3, square_direct_4, square_direct_6, square_direct_7, square_direct_8, square_direct_9, square_direct_10, square_direct_12, square_direct_13, square_direct_14, square_direct_15, square_direct_16, square_direct_17, square_direct_18,
-- 0010 multiplication with reduction and prime line not equal to 1
multiplication_with_reduction_0, multiplication_with_reduction_1, multiplication_with_reduction_2, multiplication_with_reduction_3, multiplication_with_reduction_5, multiplication_with_reduction_6, multiplication_with_reduction_7, multiplication_with_reduction_8, multiplication_with_reduction_9, multiplication_with_reduction_10, multiplication_with_reduction_11, multiplication_with_reduction_12, multiplication_with_reduction_13, multiplication_with_reduction_14, multiplication_with_reduction_16, multiplication_with_reduction_17, multiplication_with_reduction_18, multiplication_with_reduction_19, multiplication_with_reduction_20, multiplication_with_reduction_21, multiplication_with_reduction_22, multiplication_with_reduction_23, multiplication_with_reduction_24, multiplication_with_reduction_25, multiplication_with_reduction_26, multiplication_with_reduction_27, multiplication_with_reduction_28, multiplication_with_reduction_29, multiplication_with_reduction_30, multiplication_with_reduction_31, multiplication_with_reduction_32, multiplication_with_reduction_33, multiplication_with_reduction_35, multiplication_with_reduction_36, multiplication_with_reduction_37, multiplication_with_reduction_38, multiplication_with_reduction_39, multiplication_with_reduction_40, multiplication_with_reduction_41, multiplication_with_reduction_42, multiplication_with_reduction_43, multiplication_with_reduction_44, multiplication_with_reduction_45, multiplication_with_reduction_46, multiplication_with_reduction_47, multiplication_with_reduction_48, multiplication_with_reduction_49, multiplication_with_reduction_50, multiplication_with_reduction_51, multiplication_with_reduction_52, multiplication_with_reduction_53, multiplication_with_reduction_54, multiplication_with_reduction_55, multiplication_with_reduction_56, multiplication_with_reduction_57, multiplication_with_reduction_58, multiplication_with_reduction_59, multiplication_with_reduction_60, multiplication_with_reduction_61, multiplication_with_reduction_62,
-- 0010 multiplication with reduction and prime line equal to 1
multiplication_with_reduction_special_prime_0, multiplication_with_reduction_special_prime_1, multiplication_with_reduction_special_prime_3, multiplication_with_reduction_special_prime_4, multiplication_with_reduction_special_prime_5, multiplication_with_reduction_special_prime_6, multiplication_with_reduction_special_prime_7, multiplication_with_reduction_special_prime_8, multiplication_with_reduction_special_prime_10, multiplication_with_reduction_special_prime_11, multiplication_with_reduction_special_prime_12, multiplication_with_reduction_special_prime_13, multiplication_with_reduction_special_prime_14, multiplication_with_reduction_special_prime_15, multiplication_with_reduction_special_prime_16, multiplication_with_reduction_special_prime_17, multiplication_with_reduction_special_prime_18, multiplication_with_reduction_special_prime_19, multiplication_with_reduction_special_prime_20,multiplication_with_reduction_special_prime_21, multiplication_with_reduction_special_prime_22, multiplication_with_reduction_special_prime_23, multiplication_with_reduction_special_prime_25, multiplication_with_reduction_special_prime_26, multiplication_with_reduction_special_prime_27, multiplication_with_reduction_special_prime_28, multiplication_with_reduction_special_prime_29, multiplication_with_reduction_special_prime_30, multiplication_with_reduction_special_prime_31, multiplication_with_reduction_special_prime_32, multiplication_with_reduction_special_prime_33, multiplication_with_reduction_special_prime_34, multiplication_with_reduction_special_prime_35, multiplication_with_reduction_special_prime_36, multiplication_with_reduction_special_prime_37, multiplication_with_reduction_special_prime_38, multiplication_with_reduction_special_prime_39, multiplication_with_reduction_special_prime_40, multiplication_with_reduction_special_prime_41, multiplication_with_reduction_special_prime_42, multiplication_with_reduction_special_prime_43, multiplication_with_reduction_special_prime_44, multiplication_with_reduction_special_prime_45, multiplication_with_reduction_special_prime_46, multiplication_with_reduction_special_prime_47, multiplication_with_reduction_special_prime_48,
-- 0011 square with reduction and prime line not equal to 1
square_with_reduction_0, square_with_reduction_1, square_with_reduction_2, square_with_reduction_3, square_with_reduction_5, square_with_reduction_6, square_with_reduction_7, square_with_reduction_8, square_with_reduction_9, square_with_reduction_10, square_with_reduction_11, square_with_reduction_12, square_with_reduction_13, square_with_reduction_15, square_with_reduction_16, square_with_reduction_17, square_with_reduction_18, square_with_reduction_19, square_with_reduction_20, square_with_reduction_21, square_with_reduction_22, square_with_reduction_23, square_with_reduction_24, square_with_reduction_25, square_with_reduction_26, square_with_reduction_27, square_with_reduction_28, square_with_reduction_29, square_with_reduction_31, square_with_reduction_32, square_with_reduction_33, square_with_reduction_34, square_with_reduction_35, square_with_reduction_36, square_with_reduction_37, square_with_reduction_38, square_with_reduction_39, square_with_reduction_40, square_with_reduction_41, square_with_reduction_42, square_with_reduction_43, square_with_reduction_44, square_with_reduction_45, square_with_reduction_46, square_with_reduction_47, square_with_reduction_48, square_with_reduction_49, square_with_reduction_50, square_with_reduction_51, square_with_reduction_52, square_with_reduction_53,
-- 0011 square with reduction and prime line equal to 1
square_with_reduction_special_prime_0, square_with_reduction_special_prime_1, square_with_reduction_special_prime_3, square_with_reduction_special_prime_4, square_with_reduction_special_prime_5, square_with_reduction_special_prime_6, square_with_reduction_special_prime_7, square_with_reduction_special_prime_9, square_with_reduction_special_prime_10, square_with_reduction_special_prime_11, square_with_reduction_special_prime_12, square_with_reduction_special_prime_13, square_with_reduction_special_prime_14, square_with_reduction_special_prime_15, square_with_reduction_special_prime_16, square_with_reduction_special_prime_17, square_with_reduction_special_prime_18, square_with_reduction_special_prime_19, square_with_reduction_special_prime_21, square_with_reduction_special_prime_22, square_with_reduction_special_prime_23, square_with_reduction_special_prime_24, square_with_reduction_special_prime_25, square_with_reduction_special_prime_26, square_with_reduction_special_prime_27, square_with_reduction_special_prime_28, square_with_reduction_special_prime_29, square_with_reduction_special_prime_30, square_with_reduction_special_prime_31, square_with_reduction_special_prime_32, square_with_reduction_special_prime_33, square_with_reduction_special_prime_34, square_with_reduction_special_prime_35, square_with_reduction_special_prime_36, square_with_reduction_special_prime_37, square_with_reduction_special_prime_38, square_with_reduction_special_prime_39,
-- 0100 addition with no reduction
addition_subtraction_direct_0, addition_subtraction_direct_2, addition_subtraction_direct_3, addition_subtraction_direct_5, addition_subtraction_direct_6, addition_subtraction_direct_8, addition_subtraction_direct_9,
-- 0101 iterative modular reduction
iterative_modular_reduction_0, iterative_modular_reduction_1, iterative_modular_reduction_2, iterative_modular_reduction_3, iterative_modular_reduction_5, iterative_modular_reduction_6, iterative_modular_reduction_7, iterative_modular_reduction_8, iterative_modular_reduction_9, iterative_modular_reduction_10, iterative_modular_reduction_11, iterative_modular_reduction_13, iterative_modular_reduction_14, iterative_modular_reduction_15, iterative_modular_reduction_16, iterative_modular_reduction_17, iterative_modular_reduction_18, iterative_modular_reduction_19, iterative_modular_reduction_20, iterative_modular_reduction_21, iterative_modular_reduction_22, iterative_modular_reduction_24, iterative_modular_reduction_25, iterative_modular_reduction_26, iterative_modular_reduction_27, iterative_modular_reduction_28, iterative_modular_reduction_29, iterative_modular_reduction_30, iterative_modular_reduction_31, iterative_modular_reduction_32, iterative_modular_reduction_33, iterative_modular_reduction_34, iterative_modular_reduction_35, iterative_modular_reduction_36,
            
-- NOP
nop_4_stages, nop_8_stages
); 

signal actual_state, next_state : state;

signal next_sm_rotation_size : std_logic_vector(1 downto 0);
signal next_sm_circular_shift_enable : std_logic;
signal next_sel_address_a : std_logic;
signal next_sel_address_b_prime : std_logic_vector(1 downto 0);
signal next_sm_specific_mac_address_a : std_logic_vector(1 downto 0);
signal next_sm_specific_mac_address_b : std_logic_vector(1 downto 0);
signal next_sm_specific_mac_address_o : std_logic_vector(1 downto 0);
signal next_sm_specific_mac_next_address_o : std_logic_vector(1 downto 0);
signal next_mac_enable_signed_a : std_logic;
signal next_mac_enable_signed_b : std_logic;
signal next_mac_sel_load_reg_a : std_logic_vector(1 downto 0);
signal next_mac_clear_reg_b : std_logic;
signal next_mac_clear_reg_acc : std_logic;
signal next_mac_sel_shift_reg_o : std_logic;
signal next_mac_enable_update_reg_s : std_logic;
signal next_mac_sel_reg_s_reg_o_sign : std_logic;
signal next_mac_reg_s_reg_o_positive : std_logic;
signal next_sm_sign_a_mode : std_logic;
signal next_sm_mac_operation_mode : std_logic_vector(1 downto 0);
signal next_mac_enable_reg_s_mask : std_logic;
signal next_mac_subtraction_reg_a_b : std_logic;
signal next_mac_sel_multiply_two_a_b : std_logic;
signal next_mac_sel_reg_y_output : std_logic;
signal next_sm_mac_write_enable_output : std_logic;
signal next_mac_memory_double_mode : std_logic;
signal next_mac_memory_only_write_mode : std_logic;
signal next_base_address_generator_o_increment_previous_address : std_logic;
signal next_sm_free_flag : std_logic;

begin

registers_state : process(clk, rstn)
begin
    if(rstn = '0') then
        actual_state <= reset;
    elsif(rising_edge(clk)) then
        actual_state <= next_state;
    end if;
end process;

registers_state_output : process(clk)
begin
    if(rising_edge(clk)) then
        if(rstn = '0') then
            sm_free_flag <= '0';
            sm_rotation_size <= "11";
            sm_circular_shift_enable <= '0';
            sel_address_a <= '0';
            sel_address_b_prime <= "00";
            sm_specific_mac_address_a <= "00";
            sm_specific_mac_address_b <= "00";
            sm_specific_mac_address_o <= "00";
            sm_specific_mac_next_address_o <= "01";
            mac_enable_signed_a <= '0';
            mac_enable_signed_b <= '0';
            mac_sel_load_reg_a <= "11";
            mac_clear_reg_b <= '1';
            mac_clear_reg_acc <= '1';
            mac_sel_shift_reg_o <= '0';
            mac_enable_update_reg_s <= '0';
            mac_sel_reg_s_reg_o_sign <= '0';
            mac_reg_s_reg_o_positive <= '0';
            sm_sign_a_mode <= '0';
            sm_mac_operation_mode <= "10";
            mac_enable_reg_s_mask <= '0';
            mac_subtraction_reg_a_b <= '0';
            mac_sel_multiply_two_a_b <= '0';
            mac_sel_reg_y_output <= '0';
            base_address_generator_o_increment_previous_address <= '0';
            sm_mac_write_enable_output <= '0';
            mac_memory_double_mode <= '0';
            mac_memory_only_write_mode <= '0';
        else
            sm_free_flag <= next_sm_free_flag;
            sm_rotation_size <= next_sm_rotation_size;
            sm_circular_shift_enable <= next_sm_circular_shift_enable;
            sel_address_a <= next_sel_address_a;
            sel_address_b_prime <= next_sel_address_b_prime;
            sm_specific_mac_address_a <= next_sm_specific_mac_address_a;
            sm_specific_mac_address_b <= next_sm_specific_mac_address_b;
            sm_specific_mac_address_o <= next_sm_specific_mac_address_o;
            sm_specific_mac_next_address_o <= next_sm_specific_mac_next_address_o;
            mac_enable_signed_a <= next_mac_enable_signed_a;
            mac_enable_signed_b <= next_mac_enable_signed_b;
            mac_sel_load_reg_a <= next_mac_sel_load_reg_a;
            mac_clear_reg_b <= next_mac_clear_reg_b;
            mac_clear_reg_acc <= next_mac_clear_reg_acc;
            mac_sel_shift_reg_o <= next_mac_sel_shift_reg_o;
            mac_enable_update_reg_s <= next_mac_enable_update_reg_s;
            mac_sel_reg_s_reg_o_sign <= next_mac_sel_reg_s_reg_o_sign;
            mac_reg_s_reg_o_positive <= next_mac_reg_s_reg_o_positive;
            sm_sign_a_mode <= next_sm_sign_a_mode;
            sm_mac_operation_mode <= next_sm_mac_operation_mode;
            mac_enable_reg_s_mask <= next_mac_enable_reg_s_mask;
            mac_subtraction_reg_a_b <= next_mac_subtraction_reg_a_b;
            mac_sel_multiply_two_a_b <= next_mac_sel_multiply_two_a_b;
            mac_sel_reg_y_output <= next_mac_sel_reg_y_output;
            base_address_generator_o_increment_previous_address <= next_base_address_generator_o_increment_previous_address;
            sm_mac_write_enable_output <= next_sm_mac_write_enable_output;
            mac_memory_double_mode <= next_mac_memory_double_mode;
            mac_memory_only_write_mode <= next_mac_memory_only_write_mode;
        end if;
    end if;
end process;

update_output : process(actual_state, instruction_values_valid, instruction_type, operands_size)
begin
    case (actual_state) is
        when reset =>
            next_sm_free_flag <= '1';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '0';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "00";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "11";
            next_mac_clear_reg_b <= '1';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when decode_instruction =>
            next_sm_free_flag <= '1';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '0';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "00";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "11";
            next_mac_clear_reg_b <= '1';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
            if(instruction_values_valid = '1') then
                if(instruction_type = "0000") then
                    if(operands_size = "00") then
                        -- multiplication_direct_0;
                        -- -- In case of size 1
                        -- reg_a = a0_0; reg_b = b0_0; reg_acc = 0; o0_0 = reg_o; o1_0 = reg_o >> 272; Enable sign a,b; operation : a*b + acc;
                        next_sm_free_flag <= '0';
                        next_sm_rotation_size <= "11";
                        next_sm_circular_shift_enable <= '1';
                        next_sel_address_a <= '0';
                        next_sel_address_b_prime <= "00";
                        next_sm_specific_mac_address_a <= "00";
                        next_sm_specific_mac_address_b <= "00";
                        next_sm_specific_mac_address_o <= "00";
                        next_sm_specific_mac_next_address_o <= "01";
                        next_mac_enable_signed_a <= '1';
                        next_mac_enable_signed_b <= '1';
                        next_mac_sel_load_reg_a <= "00";
                        next_mac_clear_reg_b <= '0';
                        next_mac_clear_reg_acc <= '1';
                        next_mac_sel_shift_reg_o <= '0';
                        next_mac_enable_update_reg_s <= '0';
                        next_mac_sel_reg_s_reg_o_sign <= '0';
                        next_mac_reg_s_reg_o_positive <= '0';
                        next_sm_sign_a_mode <= '0';
                        next_sm_mac_operation_mode <= "10";
                        next_mac_enable_reg_s_mask <= '0';
                        next_mac_subtraction_reg_a_b <= '0';
                        next_mac_sel_multiply_two_a_b <= '0';
                        next_mac_sel_reg_y_output <= '0';
                        next_sm_mac_write_enable_output <= '1';
                        next_mac_memory_double_mode <= '1';
                        next_mac_memory_only_write_mode <= '1';
                        next_base_address_generator_o_increment_previous_address <= '0';
                    else
                        -- multiplication_direct_2;
                        -- -- Other cases
                        -- reg_a = a0_0; reg_b = b0_0; reg_acc = 0; o0_0 = reg_o; operation : a*b + acc;
                        next_sm_free_flag <= '0';
                        next_sm_rotation_size <= "11";
                        next_sm_circular_shift_enable <= '1';
                        next_sel_address_a <= '0';
                        next_sel_address_b_prime <= "00";
                        next_sm_specific_mac_address_a <= "00";
                        next_sm_specific_mac_address_b <= "00";
                        next_sm_specific_mac_address_o <= "00";
                        next_sm_specific_mac_next_address_o <= "01";
                        next_mac_enable_signed_a <= '0';
                        next_mac_enable_signed_b <= '0';
                        next_mac_sel_load_reg_a <= "00";
                        next_mac_clear_reg_b <= '0';
                        next_mac_clear_reg_acc <= '1';
                        next_mac_sel_shift_reg_o <= '0';
                        next_mac_enable_update_reg_s <= '0';
                        next_mac_sel_reg_s_reg_o_sign <= '0';
                        next_mac_reg_s_reg_o_positive <= '0';
                        next_sm_sign_a_mode <= '0';
                        next_sm_mac_operation_mode <= "10";
                        next_mac_enable_reg_s_mask <= '0';
                        next_mac_subtraction_reg_a_b <= '0';
                        next_mac_sel_multiply_two_a_b <= '0';
                        next_mac_sel_reg_y_output <= '0';
                        next_sm_mac_write_enable_output <= '1';
                        next_mac_memory_double_mode <= '0';
                        next_mac_memory_only_write_mode <= '0';
                        next_base_address_generator_o_increment_previous_address <= '0';
                    end if;
                elsif(instruction_type = "0001") then
                    if(operands_size = "00") then
                        -- square_direct_0;
                        -- -- In case of size 1
                        -- reg_a = a0_0; reg_b = a0_0; reg_acc = 0; o0_0 = reg_o; o1_0 = reg_o >> 272; Enable sign a,b; operation : a*b + acc;
                        next_sm_free_flag <= '0';
                        next_sm_rotation_size <= "11";
                        next_sm_circular_shift_enable <= '1';
                        next_sel_address_a <= '0';
                        next_sel_address_b_prime <= "00";
                        next_sm_specific_mac_address_a <= "00";
                        next_sm_specific_mac_address_b <= "00";
                        next_sm_specific_mac_address_o <= "00";
                        next_sm_specific_mac_next_address_o <= "01";
                        next_mac_enable_signed_a <= '1';
                        next_mac_enable_signed_b <= '1';
                        next_mac_sel_load_reg_a <= "00";
                        next_mac_clear_reg_b <= '0';
                        next_mac_clear_reg_acc <= '1';
                        next_mac_sel_shift_reg_o <= '0';
                        next_mac_enable_update_reg_s <= '0';
                        next_mac_sel_reg_s_reg_o_sign <= '0';
                        next_mac_reg_s_reg_o_positive <= '0';
                        next_sm_sign_a_mode <= '0';
                        next_sm_mac_operation_mode <= "10";
                        next_mac_enable_reg_s_mask <= '0';
                        next_mac_subtraction_reg_a_b <= '0';
                        next_mac_sel_multiply_two_a_b <= '0';
                        next_mac_sel_reg_y_output <= '0';
                        next_sm_mac_write_enable_output <= '1';
                        next_mac_memory_double_mode <= '1';
                        next_mac_memory_only_write_mode <= '1';
                        next_base_address_generator_o_increment_previous_address <= '0';
                    else
                        -- square_direct_2;
                        -- -- In case of sizes 2, 3, 4
                        -- reg_a = a0_0; reg_b = a0_0; reg_acc = 0; o0_0 = reg_o; operation : a*b + acc;
                        next_sm_free_flag <= '0';
                        next_sm_rotation_size <= "11";
                        next_sm_circular_shift_enable <= '1';
                        next_sel_address_a <= '0';
                        next_sel_address_b_prime <= "00";
                        next_sm_specific_mac_address_a <= "00";
                        next_sm_specific_mac_address_b <= "00";
                        next_sm_specific_mac_address_o <= "00";
                        next_sm_specific_mac_next_address_o <= "01";
                        next_mac_enable_signed_a <= '0';
                        next_mac_enable_signed_b <= '0';
                        next_mac_sel_load_reg_a <= "00";
                        next_mac_clear_reg_b <= '0';
                        next_mac_clear_reg_acc <= '1';
                        next_mac_sel_shift_reg_o <= '0';
                        next_mac_enable_update_reg_s <= '0';
                        next_mac_sel_reg_s_reg_o_sign <= '0';
                        next_mac_reg_s_reg_o_positive <= '0';
                        next_sm_sign_a_mode <= '0';
                        next_sm_mac_operation_mode <= "10";
                        next_mac_enable_reg_s_mask <= '0';
                        next_mac_subtraction_reg_a_b <= '0';
                        next_mac_sel_multiply_two_a_b <= '0';
                        next_mac_sel_reg_y_output <= '0';
                        next_sm_mac_write_enable_output <= '1';
                        next_mac_memory_double_mode <= '0';
                        next_mac_memory_only_write_mode <= '0';
                        next_base_address_generator_o_increment_previous_address <= '0';
                    end if;
                elsif(instruction_type = "0010") then
                    if(prime_line_equal_one = '1') then
                        if(operands_size = "00") then
                            -- multiplication_with_reduction_special_prime_0;
                            -- -- In case of size 1
                            -- reg_a = a0_0; reg_b = b0_0; reg_acc = 0; Enable sign a,b; operation : a*b + acc;
                            next_sm_free_flag <= '0';
                            next_sm_rotation_size <= "11";
                            next_sm_circular_shift_enable <= '1';
                            next_sel_address_a <= '0';
                            next_sel_address_b_prime <= "00";
                            next_sm_specific_mac_address_a <= "00";
                            next_sm_specific_mac_address_b <= "00";
                            next_sm_specific_mac_address_o <= "00";
                            next_sm_specific_mac_next_address_o <= "01";
                            next_mac_enable_signed_a <= '0';
                            next_mac_enable_signed_b <= '0';
                            next_mac_sel_load_reg_a <= "00";
                            next_mac_clear_reg_b <= '0';
                            next_mac_clear_reg_acc <= '1';
                            next_mac_sel_shift_reg_o <= '0';
                            next_mac_enable_update_reg_s <= '0';
                            next_mac_sel_reg_s_reg_o_sign <= '0';
                            next_mac_reg_s_reg_o_positive <= '0';
                            next_sm_sign_a_mode <= '0';
                            next_sm_mac_operation_mode <= "10";
                            next_mac_enable_reg_s_mask <= '0';
                            next_mac_subtraction_reg_a_b <= '0';
                            next_mac_sel_multiply_two_a_b <= '0';
                            next_mac_sel_reg_y_output <= '0';
                            next_sm_mac_write_enable_output <= '0';
                            next_mac_memory_double_mode <= '0';
                            next_mac_memory_only_write_mode <= '0';
                            next_base_address_generator_o_increment_previous_address <= '0';
                        else
                            -- multiplication_with_reduction_special_prime_3;
                            -- -- In case of sizes 2, 3, 4
                            -- reg_a = a0_0; reg_b = b0_0; reg_acc = 0; o0_0 = reg_o; operation : a*b + acc;
                            next_sm_free_flag <= '0';
                            next_sm_rotation_size <= "11";
                            next_sm_circular_shift_enable <= '1';
                            next_sel_address_a <= '0';
                            next_sel_address_b_prime <= "00";
                            next_sm_specific_mac_address_a <= "00";
                            next_sm_specific_mac_address_b <= "00";
                            next_sm_specific_mac_address_o <= "00";
                            next_sm_specific_mac_next_address_o <= "01";
                            next_mac_enable_signed_a <= '0';
                            next_mac_enable_signed_b <= '0';
                            next_mac_sel_load_reg_a <= "00";
                            next_mac_clear_reg_b <= '0';
                            next_mac_clear_reg_acc <= '1';
                            next_mac_sel_shift_reg_o <= '0';
                            next_mac_enable_update_reg_s <= '0';
                            next_mac_sel_reg_s_reg_o_sign <= '0';
                            next_mac_reg_s_reg_o_positive <= '0';
                            next_sm_sign_a_mode <= '0';
                            next_sm_mac_operation_mode <= "10";
                            next_mac_enable_reg_s_mask <= '0';
                            next_mac_subtraction_reg_a_b <= '0';
                            next_mac_sel_multiply_two_a_b <= '0';
                            next_mac_sel_reg_y_output <= '0';
                            next_sm_mac_write_enable_output <= '1';
                            next_mac_memory_double_mode <= '0';
                            next_mac_memory_only_write_mode <= '0';
                            next_base_address_generator_o_increment_previous_address <= '0';
                        end if;
                    else
                        if(operands_size = "00") then
                            -- multiplication_with_reduction_0
                            -- -- In case of size 1
                            -- reg_a = a0_0; reg_b = b0_0; reg_acc = 0; Enable sign a,b; operation : a*b + acc;
                            next_sm_free_flag <= '0';
                            next_sm_rotation_size <= "11";
                            next_sm_circular_shift_enable <= '1';
                            next_sel_address_a <= '0';
                            next_sel_address_b_prime <= "00";
                            next_sm_specific_mac_address_a <= "00";
                            next_sm_specific_mac_address_b <= "00";
                            next_sm_specific_mac_address_o <= "00";
                            next_sm_specific_mac_next_address_o <= "01";
                            next_mac_enable_signed_a <= '1';
                            next_mac_enable_signed_b <= '1';
                            next_mac_sel_load_reg_a <= "00";
                            next_mac_clear_reg_b <= '0';
                            next_mac_clear_reg_acc <= '1';
                            next_mac_sel_shift_reg_o <= '0';
                            next_mac_enable_update_reg_s <= '0';
                            next_mac_sel_reg_s_reg_o_sign <= '0';
                            next_mac_reg_s_reg_o_positive <= '0';
                            next_sm_sign_a_mode <= '0';
                            next_sm_mac_operation_mode <= "10";
                            next_mac_enable_reg_s_mask <= '0';
                            next_mac_subtraction_reg_a_b <= '0';
                            next_mac_sel_multiply_two_a_b <= '0';
                            next_mac_sel_reg_y_output <= '0';
                            next_sm_mac_write_enable_output <= '0';
                            next_mac_memory_double_mode <= '0';
                            next_mac_memory_only_write_mode <= '0';
                            next_base_address_generator_o_increment_previous_address <= '0';
                        else
                            -- multiplication_with_reduction_5
                            -- -- In case of sizes 2, 3, 4
                            -- reg_a = a0_0; reg_b = b0_0; reg_acc = 0; operation : a*b + acc;
                            next_sm_free_flag <= '0';
                            next_sm_rotation_size <= "11";
                            next_sm_circular_shift_enable <= '1';
                            next_sel_address_a <= '0';
                            next_sel_address_b_prime <= "00";
                            next_sm_specific_mac_address_a <= "00";
                            next_sm_specific_mac_address_b <= "00";
                            next_sm_specific_mac_address_o <= "00";
                            next_sm_specific_mac_next_address_o <= "01";
                            next_mac_enable_signed_a <= '0';
                            next_mac_enable_signed_b <= '0';
                            next_mac_sel_load_reg_a <= "00";
                            next_mac_clear_reg_b <= '0';
                            next_mac_clear_reg_acc <= '1';
                            next_mac_sel_shift_reg_o <= '0';
                            next_mac_enable_update_reg_s <= '0';
                            next_mac_sel_reg_s_reg_o_sign <= '0';
                            next_mac_reg_s_reg_o_positive <= '0';
                            next_sm_sign_a_mode <= '0';
                            next_sm_mac_operation_mode <= "10";
                            next_mac_enable_reg_s_mask <= '0';
                            next_mac_subtraction_reg_a_b <= '0';
                            next_mac_sel_multiply_two_a_b <= '0';
                            next_mac_sel_reg_y_output <= '0';
                            next_sm_mac_write_enable_output <= '0';
                            next_mac_memory_double_mode <= '0';
                            next_mac_memory_only_write_mode <= '0';
                            next_base_address_generator_o_increment_previous_address <= '0';
                        end if;
                    end if;
                elsif(instruction_type = "0011") then
                    if(prime_line_equal_one = '1') then
                        if(operands_size = "00") then
                            -- square_with_reduction_special_prime_0
                            -- -- In case of size 1
                            -- reg_a = a0_0; reg_b = a0_0; reg_acc = 0; Enable sign a,b; operation : a*b + acc;
                            next_sm_free_flag <= '0';
                            next_sm_rotation_size <= "11";
                            next_sm_circular_shift_enable <= '1';
                            next_sel_address_a <= '0';
                            next_sel_address_b_prime <= "00";
                            next_sm_specific_mac_address_a <= "00";
                            next_sm_specific_mac_address_b <= "00";
                            next_sm_specific_mac_address_o <= "00";
                            next_sm_specific_mac_next_address_o <= "01";
                            next_mac_enable_signed_a <= '1';
                            next_mac_enable_signed_b <= '1';
                            next_mac_sel_load_reg_a <= "00";
                            next_mac_clear_reg_b <= '0';
                            next_mac_clear_reg_acc <= '1';
                            next_mac_sel_shift_reg_o <= '0';
                            next_mac_enable_update_reg_s <= '0';
                            next_mac_sel_reg_s_reg_o_sign <= '0';
                            next_mac_reg_s_reg_o_positive <= '0';
                            next_sm_sign_a_mode <= '0';
                            next_sm_mac_operation_mode <= "10";
                            next_mac_enable_reg_s_mask <= '0';
                            next_mac_subtraction_reg_a_b <= '0';
                            next_mac_sel_multiply_two_a_b <= '0';
                            next_mac_sel_reg_y_output <= '0';
                            next_sm_mac_write_enable_output <= '0';
                            next_mac_memory_double_mode <= '0';
                            next_mac_memory_only_write_mode <= '0';
                            next_base_address_generator_o_increment_previous_address <= '0';
                        else
                            -- square_with_reduction_special_prime_3
                            -- -- In case of size 2, 3, 4
                            -- reg_a = a0_0; reg_b = a0_0; reg_acc = 0; o0_0 = reg_o; operation : a*b + acc;
                            next_sm_free_flag <= '0';
                            next_sm_rotation_size <= "11";
                            next_sm_circular_shift_enable <= '1';
                            next_sel_address_a <= '0';
                            next_sel_address_b_prime <= "00";
                            next_sm_specific_mac_address_a <= "00";
                            next_sm_specific_mac_address_b <= "00";
                            next_sm_specific_mac_address_o <= "00";
                            next_sm_specific_mac_next_address_o <= "01";
                            next_mac_enable_signed_a <= '0';
                            next_mac_enable_signed_b <= '0';
                            next_mac_sel_load_reg_a <= "00";
                            next_mac_clear_reg_b <= '0';
                            next_mac_clear_reg_acc <= '1';
                            next_mac_sel_shift_reg_o <= '0';
                            next_mac_enable_update_reg_s <= '0';
                            next_mac_sel_reg_s_reg_o_sign <= '0';
                            next_mac_reg_s_reg_o_positive <= '0';
                            next_sm_sign_a_mode <= '0';
                            next_sm_mac_operation_mode <= "10";
                            next_mac_enable_reg_s_mask <= '0';
                            next_mac_subtraction_reg_a_b <= '0';
                            next_mac_sel_multiply_two_a_b <= '0';
                            next_mac_sel_reg_y_output <= '0';
                            next_sm_mac_write_enable_output <= '1';
                            next_mac_memory_double_mode <= '0';
                            next_mac_memory_only_write_mode <= '0';
                            next_base_address_generator_o_increment_previous_address <= '0';
                        end if;
                    else
                        if(operands_size = "00") then
                            -- square_with_reduction_0
                            -- -- In case of size 1
                            -- reg_a = a0_0; reg_b = a0_0; reg_acc = 0; Enable sign a,b; operation : a*b + acc;
                            next_sm_free_flag <= '0';
                            next_sm_rotation_size <= "11";
                            next_sm_circular_shift_enable <= '1';
                            next_sel_address_a <= '0';
                            next_sel_address_b_prime <= "00";
                            next_sm_specific_mac_address_a <= "00";
                            next_sm_specific_mac_address_b <= "00";
                            next_sm_specific_mac_address_o <= "00";
                            next_sm_specific_mac_next_address_o <= "01";
                            next_mac_enable_signed_a <= '1';
                            next_mac_enable_signed_b <= '1';
                            next_mac_sel_load_reg_a <= "00";
                            next_mac_clear_reg_b <= '0';
                            next_mac_clear_reg_acc <= '1';
                            next_mac_sel_shift_reg_o <= '0';
                            next_mac_enable_update_reg_s <= '0';
                            next_mac_sel_reg_s_reg_o_sign <= '0';
                            next_mac_reg_s_reg_o_positive <= '0';
                            next_sm_sign_a_mode <= '0';
                            next_sm_mac_operation_mode <= "10";
                            next_mac_enable_reg_s_mask <= '0';
                            next_mac_subtraction_reg_a_b <= '0';
                            next_mac_sel_multiply_two_a_b <= '0';
                            next_mac_sel_reg_y_output <= '0';
                            next_sm_mac_write_enable_output <= '0';
                            next_mac_memory_double_mode <= '0';
                            next_mac_memory_only_write_mode <= '0';
                            next_base_address_generator_o_increment_previous_address <= '0';
                        else
                            -- square_with_reduction_5
                            -- -- In case of 2, 3, 4
                            -- reg_a = a0_0; reg_b = a0_0; reg_acc = 0; operation : a*b + acc;
                            next_sm_free_flag <= '0';
                            next_sm_rotation_size <= "11";
                            next_sm_circular_shift_enable <= '1';
                            next_sel_address_a <= '0';
                            next_sel_address_b_prime <= "00";
                            next_sm_specific_mac_address_a <= "00";
                            next_sm_specific_mac_address_b <= "00";
                            next_sm_specific_mac_address_o <= "00";
                            next_sm_specific_mac_next_address_o <= "01";
                            next_mac_enable_signed_a <= '0';
                            next_mac_enable_signed_b <= '0';
                            next_mac_sel_load_reg_a <= "00";
                            next_mac_clear_reg_b <= '0';
                            next_mac_clear_reg_acc <= '1';
                            next_mac_sel_shift_reg_o <= '0';
                            next_mac_enable_update_reg_s <= '0';
                            next_mac_sel_reg_s_reg_o_sign <= '0';
                            next_mac_reg_s_reg_o_positive <= '0';
                            next_sm_sign_a_mode <= '0';
                            next_sm_mac_operation_mode <= "10";
                            next_mac_enable_reg_s_mask <= '0';
                            next_mac_subtraction_reg_a_b <= '0';
                            next_mac_sel_multiply_two_a_b <= '0';
                            next_mac_sel_reg_y_output <= '0';
                            next_sm_mac_write_enable_output <= '0';
                            next_mac_memory_double_mode <= '0';
                            next_mac_memory_only_write_mode <= '0';
                            next_base_address_generator_o_increment_previous_address <= '0';
                        end if;
                    end if;
                elsif(instruction_type = "0100") then
                    if(operands_size = "00") then
                        -- addition_subtraction_direct_0
                        -- -- In case of size 1
                        -- reg_a = a0_0; reg_b = b0_0; reg_acc = 0; o0_0 = reg_o; Enable sign a,b; operation : b +/- a + acc;
                        next_sm_free_flag <= '0';
                        next_sm_rotation_size <= "10";
                        next_sm_circular_shift_enable <= '1';
                        next_sel_address_a <= '0';
                        next_sel_address_b_prime <= "00";
                        next_sm_specific_mac_address_a <= "00";
                        next_sm_specific_mac_address_b <= "00";
                        next_sm_specific_mac_address_o <= "00";
                        next_sm_specific_mac_next_address_o <= "01";
                        next_mac_enable_signed_a <= '1';
                        next_mac_enable_signed_b <= '1';
                        next_mac_sel_load_reg_a <= "00";
                        next_mac_clear_reg_b <= '0';
                        next_mac_clear_reg_acc <= '1';
                        next_mac_sel_shift_reg_o <= '0';
                        next_mac_enable_update_reg_s <= '0';
                        next_mac_sel_reg_s_reg_o_sign <= '0';
                        next_mac_reg_s_reg_o_positive <= '0';
                        next_sm_sign_a_mode <= '1';
                        next_sm_mac_operation_mode(1) <= '0';
                        next_sm_mac_operation_mode(0) <= '0';
                        next_mac_enable_reg_s_mask <= '0';
                        next_mac_subtraction_reg_a_b <= '0';
                        next_mac_sel_multiply_two_a_b <= '0';
                        next_mac_sel_reg_y_output <= '0';
                        next_sm_mac_write_enable_output <= '1';
                        next_mac_memory_double_mode <= '0';
                        next_mac_memory_only_write_mode <= '0';
                        next_base_address_generator_o_increment_previous_address <= '0';
                    else
                        -- addition_subtraction_direct_2
                        -- -- In case of size 2, 3, 4
                        -- reg_a = a0_0; reg_b = b0_0; reg_acc = 0; o0_0 = reg_o; operation : b +/- a + acc;
                        next_sm_free_flag <= '0';
                        next_sm_rotation_size <= "10";
                        next_sm_circular_shift_enable <= '1';
                        next_sel_address_a <= '0';
                        next_sel_address_b_prime <= "00";
                        next_sm_specific_mac_address_a <= "00";
                        next_sm_specific_mac_address_b <= "00";
                        next_sm_specific_mac_address_o <= "00";
                        next_sm_specific_mac_next_address_o <= "01";
                        next_mac_enable_signed_a <= '0';
                        next_mac_enable_signed_b <= '0';
                        next_mac_sel_load_reg_a <= "00";
                        next_mac_clear_reg_b <= '0';
                        next_mac_clear_reg_acc <= '1';
                        next_mac_sel_shift_reg_o <= '0';
                        next_mac_enable_update_reg_s <= '0';
                        next_mac_sel_reg_s_reg_o_sign <= '0';
                        next_mac_reg_s_reg_o_positive <= '0';
                        next_sm_sign_a_mode <= '1';
                        next_sm_mac_operation_mode(1) <= '0';
                        next_sm_mac_operation_mode(0) <= '0';
                        next_mac_enable_reg_s_mask <= '0';
                        next_mac_subtraction_reg_a_b <= '0';
                        next_mac_sel_multiply_two_a_b <= '0';
                        next_mac_sel_reg_y_output <= '0';
                        next_sm_mac_write_enable_output <= '1';
                        next_mac_memory_double_mode <= '0';
                        next_mac_memory_only_write_mode <= '0';
                        next_base_address_generator_o_increment_previous_address <= '0';
                    end if;
                elsif(instruction_type = "0101") then
                    if(operands_size = "00") then
                        -- iterative_modular_reduction_0
                        -- reg_a = a0_0; reg_b = 0; reg_acc = 0; Enable sign a,b; operation : b + a + acc;
                        next_sm_free_flag <= '0';
                        next_sm_rotation_size <= "10";
                        next_sm_circular_shift_enable <= '1';
                        next_sel_address_a <= '0';
                        next_sel_address_b_prime <= "10";
                        next_sm_specific_mac_address_a <= "00";
                        next_sm_specific_mac_address_b <= "00";
                        next_sm_specific_mac_address_o <= "00";
                        next_sm_specific_mac_next_address_o <= "01";
                        next_mac_enable_signed_a <= '1';
                        next_mac_enable_signed_b <= '1';
                        next_mac_sel_load_reg_a <= "00";
                        next_mac_clear_reg_b <= '1';
                        next_mac_clear_reg_acc <= '1';
                        next_mac_sel_shift_reg_o <= '0';
                        next_mac_enable_update_reg_s <= '0';
                        next_mac_sel_reg_s_reg_o_sign <= '0';
                        next_mac_reg_s_reg_o_positive <= '0';
                        next_sm_sign_a_mode <= '0';
                        next_sm_mac_operation_mode <= "01";
                        next_mac_enable_reg_s_mask <= '0';
                        next_mac_subtraction_reg_a_b <= '0';
                        next_mac_sel_multiply_two_a_b <= '0';
                        next_mac_sel_reg_y_output <= '0';
                        next_sm_mac_write_enable_output <= '0';
                        next_mac_memory_double_mode <= '0';
                        next_mac_memory_only_write_mode <= '0';
                        next_base_address_generator_o_increment_previous_address <= '0';
                    elsif(operands_size = "01") then
                        -- iterative_modular_reduction_5
                        -- reg_a = a1_0; reg_b = 0; reg_acc = 0; Enable sign a,b; operation : b + a + acc;
                        next_sm_free_flag <= '0';
                        next_sm_rotation_size <= "10";
                        next_sm_circular_shift_enable <= '1';
                        next_sel_address_a <= '0';
                        next_sel_address_b_prime <= "10";
                        next_sm_specific_mac_address_a <= "01";
                        next_sm_specific_mac_address_b <= "00";
                        next_sm_specific_mac_address_o <= "00";
                        next_sm_specific_mac_next_address_o <= "01";
                        next_mac_enable_signed_a <= '1';
                        next_mac_enable_signed_b <= '1';
                        next_mac_sel_load_reg_a <= "00";
                        next_mac_clear_reg_b <= '1';
                        next_mac_clear_reg_acc <= '1';
                        next_mac_sel_shift_reg_o <= '0';
                        next_mac_enable_update_reg_s <= '0';
                        next_mac_sel_reg_s_reg_o_sign <= '0';
                        next_mac_reg_s_reg_o_positive <= '0';
                        next_sm_sign_a_mode <= '0';
                        next_sm_mac_operation_mode <= "01";
                        next_mac_enable_reg_s_mask <= '0';
                        next_mac_subtraction_reg_a_b <= '0';
                        next_mac_sel_multiply_two_a_b <= '0';
                        next_mac_sel_reg_y_output <= '0';
                        next_sm_mac_write_enable_output <= '0';
                        next_mac_memory_double_mode <= '0';
                        next_mac_memory_only_write_mode <= '0';
                        next_base_address_generator_o_increment_previous_address <= '0';
                    elsif(operands_size = "10") then
                        -- iterative_modular_reduction_13
                        -- reg_a = a2_0; reg_b = 0; reg_acc = 0; Enable sign a,b; operation : b + a + acc;
                        next_sm_free_flag <= '0';
                        next_sm_rotation_size <= "10";
                        next_sm_circular_shift_enable <= '1';
                        next_sel_address_a <= '0';
                        next_sel_address_b_prime <= "10";
                        next_sm_specific_mac_address_a <= "10";
                        next_sm_specific_mac_address_b <= "10";
                        next_sm_specific_mac_address_o <= "10";
                        next_sm_specific_mac_next_address_o <= "11";
                        next_mac_enable_signed_a <= '1';
                        next_mac_enable_signed_b <= '1';
                        next_mac_sel_load_reg_a <= "00";
                        next_mac_clear_reg_b <= '1';
                        next_mac_clear_reg_acc <= '1';
                        next_mac_sel_shift_reg_o <= '0';
                        next_mac_enable_update_reg_s <= '0';
                        next_mac_sel_reg_s_reg_o_sign <= '0';
                        next_mac_reg_s_reg_o_positive <= '0';
                        next_sm_sign_a_mode <= '0';
                        next_sm_mac_operation_mode <= "01";
                        next_mac_enable_reg_s_mask <= '0';
                        next_mac_subtraction_reg_a_b <= '0';
                        next_mac_sel_multiply_two_a_b <= '0';
                        next_mac_sel_reg_y_output <= '0';
                        next_sm_mac_write_enable_output <= '0';
                        next_mac_memory_double_mode <= '0';
                        next_mac_memory_only_write_mode <= '0';
                        next_base_address_generator_o_increment_previous_address <= '0';
                    else
                        -- iterative_modular_reduction_24
                        -- reg_a = a3_0; reg_b = 0; reg_acc = 0; Enable sign a,b; operation : b + a + acc;
                        next_sm_free_flag <= '0';
                        next_sm_rotation_size <= "10";
                        next_sm_circular_shift_enable <= '1';
                        next_sel_address_a <= '0';
                        next_sel_address_b_prime <= "10";
                        next_sm_specific_mac_address_a <= "11";
                        next_sm_specific_mac_address_b <= "11";
                        next_sm_specific_mac_address_o <= "11";
                        next_sm_specific_mac_next_address_o <= "00";
                        next_mac_enable_signed_a <= '1';
                        next_mac_enable_signed_b <= '1';
                        next_mac_sel_load_reg_a <= "00";
                        next_mac_clear_reg_b <= '1';
                        next_mac_clear_reg_acc <= '1';
                        next_mac_sel_shift_reg_o <= '0';
                        next_mac_enable_update_reg_s <= '0';
                        next_mac_sel_reg_s_reg_o_sign <= '0';
                        next_mac_reg_s_reg_o_positive <= '0';
                        next_sm_sign_a_mode <= '0';
                        next_sm_mac_operation_mode <= "01";
                        next_mac_enable_reg_s_mask <= '0';
                        next_mac_subtraction_reg_a_b <= '0';
                        next_mac_sel_multiply_two_a_b <= '0';
                        next_mac_sel_reg_y_output <= '0';
                        next_sm_mac_write_enable_output <= '0';
                        next_mac_memory_double_mode <= '0';
                        next_mac_memory_only_write_mode <= '0';
                        next_base_address_generator_o_increment_previous_address <= '0';
                    end if;
                end if;
                
                
                if(instruction_type = "0000") then
                    next_sm_rotation_size <= "11";
                elsif(instruction_type = "0001") then
                    next_sm_rotation_size <= "11";
                elsif(instruction_type = "0010") then
                    next_sm_rotation_size <= "11";
                elsif(instruction_type = "0011") then
                    next_sm_rotation_size <= "11";
                elsif(instruction_type = "0100") then
                    next_sm_rotation_size <= "10";
                elsif(instruction_type = "0101") then
                    next_sm_rotation_size <= "10";
                elsif(instruction_type = "0110") then
                    next_sm_rotation_size <= "00";
                end if;
            end if;
        when multiplication_direct_0 =>
        -- -- In case of size 1
        -- reg_a = a0_0; reg_b = b0_0; reg_acc = 0; o0_0 = reg_o; o1_0 = reg_o >> 272; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "00";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_2 =>
         -- -- Other cases
        -- reg_a = a0_0; reg_b = b0_0; reg_acc = 0; o0_0 = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "00";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_3 =>
        -- -- In case of size 2
        -- reg_a = a1_0; reg_b = b0_0; reg_acc = reg_o >> 272; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "01";
            next_sm_specific_mac_address_b <= "00";
            next_sm_specific_mac_address_o <= "01";
            next_sm_specific_mac_next_address_o <= "10";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_4 =>
        -- reg_a = a0_0; reg_b = b1_0; reg_acc = reg_o; o1_0 = reg_o; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "01";
            next_sm_specific_mac_address_o <= "01";
            next_sm_specific_mac_next_address_o <= "10";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_5 =>
            -- reg_a = a1_0; reg_b = b1_0; reg_acc = reg_o >> 272; o2_0 = reg_o; o3_0 = reg_o >> 272; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "01";
            next_sm_specific_mac_address_b <= "01";
            next_sm_specific_mac_address_o <= "10";
            next_sm_specific_mac_next_address_o <= "11";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_7 =>
        -- -- In case of size 3, 4           
        -- reg_a = a1_0; reg_b = b0_0; reg_acc = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "01";
            next_sm_specific_mac_address_b <= "00";
            next_sm_specific_mac_address_o <= "01";
            next_sm_specific_mac_next_address_o <= "10";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_8 =>
        -- reg_a = a0_0; reg_b = b1_0; reg_acc = reg_o; o1_0 = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "01";
            next_sm_specific_mac_address_o <= "01";
            next_sm_specific_mac_next_address_o <= "10";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_9 =>
            -- reg_a = a1_0; reg_b = b1_0; reg_acc = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "01";
            next_sm_specific_mac_address_b <= "01";
            next_sm_specific_mac_address_o <= "10";
            next_sm_specific_mac_next_address_o <= "11";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_10 =>
        -- -- In case of size 3
        -- reg_a = a0_0; reg_b = b2_0; reg_acc = reg_o; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "10";
            next_sm_specific_mac_address_o <= "10";
            next_sm_specific_mac_next_address_o <= "11";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_11 =>
        -- reg_a = a2_0; reg_b = b0_0; reg_acc = reg_o; o2_0 = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "10";
            next_sm_specific_mac_address_b <= "00";
            next_sm_specific_mac_address_o <= "10";
            next_sm_specific_mac_next_address_o <= "11";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_12 =>
            -- reg_a = a2_0; reg_b = b1_0; reg_acc = reg_o >> 272; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "10";
            next_sm_specific_mac_address_b <= "01";
            next_sm_specific_mac_address_o <= "11";
            next_sm_specific_mac_next_address_o <= "00";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_13 =>
            -- reg_a = a1_0; reg_b = b2_0; reg_acc = reg_o; o3_0 = reg_o; Enable sign b; operation : a*b + acc; Increment o3_0 base address
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "01";
            next_sm_specific_mac_address_b <= "10";
            next_sm_specific_mac_address_o <= "11";
            next_sm_specific_mac_next_address_o <= "00";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '1';
        when multiplication_direct_14 =>
        -- reg_a = a2_0; reg_b = b2_0; reg_acc = reg_o >> 272; o4_0 = reg_o; o5_0 = reg_o >> 272; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "10";
            next_sm_specific_mac_address_b <= "10";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_16 =>
        -- -- In case of size 4
        -- reg_a = a0_0; reg_b = b2_0; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "10";
            next_sm_specific_mac_address_o <= "10";
            next_sm_specific_mac_next_address_o <= "11";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_17 =>
        -- reg_a = a2_0; reg_b = b0_0; reg_acc = reg_o; o2_0 = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "10";
            next_sm_specific_mac_address_b <= "00";
            next_sm_specific_mac_address_o <= "10";
            next_sm_specific_mac_next_address_o <= "11";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_18 =>
            -- reg_a = a2_0; reg_b = b1_0; reg_acc = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "10";
            next_sm_specific_mac_address_b <= "01";
            next_sm_specific_mac_address_o <= "11";
            next_sm_specific_mac_next_address_o <= "00";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_19 =>
            -- reg_a = a1_0; reg_b = b2_0; reg_acc = reg_o; operation : a*b + acc; 
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "01";
            next_sm_specific_mac_address_b <= "10";
            next_sm_specific_mac_address_o <= "11";
            next_sm_specific_mac_next_address_o <= "00";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_20 =>
        -- reg_a = a3_0; reg_b = b0_0; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "11";
            next_sm_specific_mac_address_b <= "00";
            next_sm_specific_mac_address_o <= "11";
            next_sm_specific_mac_next_address_o <= "00";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_21 =>
        -- reg_a = a0_0; reg_b = b3_0; reg_acc = reg_o; o3_0 = reg_o; Enable sign b; operation : a*b + acc; Increment o3_0 base address
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "11";
            next_sm_specific_mac_address_o <= "11";
            next_sm_specific_mac_next_address_o <= "00";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '1';
        when multiplication_direct_22 =>
            -- reg_a = a2_0; reg_b = b2_0; reg_acc = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "10";
            next_sm_specific_mac_address_b <= "10";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_23 =>
            -- reg_a = a3_0; reg_b = b1_0; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "11";
            next_sm_specific_mac_address_b <= "01";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_24 =>
            -- reg_a = a1_0; reg_b = b3_0; reg_acc = reg_o; o4_0 = reg_o; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "01";
            next_sm_specific_mac_address_b <= "11";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_25 =>
            -- reg_a = a3_0; reg_b = b2_0; reg_acc = reg_o >> 272; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "11";
            next_sm_specific_mac_address_b <= "10";
            next_sm_specific_mac_address_o <= "01";
            next_sm_specific_mac_next_address_o <= "10";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_26 =>
            -- reg_a = a2_0; reg_b = b3_0; reg_acc = reg_o; o5_0 = reg_o; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "10";
            next_sm_specific_mac_address_b <= "11";
            next_sm_specific_mac_address_o <= "01";
            next_sm_specific_mac_next_address_o <= "10";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_direct_27 =>
            -- reg_a = a3_0; reg_b = b3_0; reg_acc = reg_o >> 272; o6_0 = reg_o; o7_0 = reg_o >> 272; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "11";
            next_sm_specific_mac_address_b <= "11";
            next_sm_specific_mac_address_o <= "10";
            next_sm_specific_mac_next_address_o <= "11";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_0 => 
            -- -- In case of size 1
            -- reg_a = a0_0; reg_b = a0_0; reg_acc = 0; o0_0 = reg_o; o1_0 = reg_o >> 272; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "00";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_2 => 
            -- -- In case of sizes 2, 3, 4
            -- reg_a = a0_0; reg_b = a0_0; reg_acc = 0; o0_0 = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "00";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_3 => 
            -- -- In case of size 2
            -- reg_a = a1_0; reg_b = a0_0; reg_acc = reg_o >> 272; o1_0 = reg_o; Enable sign a; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "01";
            next_sm_specific_mac_address_b <= "00";
            next_sm_specific_mac_address_o <= "01";
            next_sm_specific_mac_next_address_o <= "10";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_4 => 
            -- reg_a = a1_0; reg_b = a1_0; reg_acc = reg_o >> 272; o2_0 = reg_o; o3_0 = reg_o >> 272; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "01";
            next_sm_specific_mac_address_b <= "01";
            next_sm_specific_mac_address_o <= "10";
            next_sm_specific_mac_next_address_o <= "11";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_6 => 
            -- -- In case of sizes 3, 4
            -- reg_a = a1_0; reg_b = a0_0; reg_acc = reg_o >> 272; o1_0 = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "01";
            next_sm_specific_mac_address_b <= "00";
            next_sm_specific_mac_address_o <= "01";
            next_sm_specific_mac_next_address_o <= "10";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_7 =>
            -- reg_a = a1_0; reg_b = a1_0; reg_acc = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "01";
            next_sm_specific_mac_address_b <= "01";
            next_sm_specific_mac_address_o <= "10";
            next_sm_specific_mac_next_address_o <= "11";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_8 =>
            -- -- In case of size 3
            -- reg_a = a0_0; reg_b = a2_0; reg_acc = reg_o; o2_0 = reg_o; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "10";
            next_sm_specific_mac_address_o <= "10";
            next_sm_specific_mac_next_address_o <= "11";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_9 =>
            -- reg_a = a2_0; reg_b = a1_0; reg_acc = reg_o >> 272; o3_0 = reg_o; Enable sign a; operation : 2*a*b + acc; Increment o3_0 base address
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "10";
            next_sm_specific_mac_address_b <= "01";
            next_sm_specific_mac_address_o <= "11";
            next_sm_specific_mac_next_address_o <= "00";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '1';
        when square_direct_10 =>
            -- reg_a = a2_0; reg_b = a2_0; reg_acc = reg_o >> 272; o4_0 = reg_o; o5_0 = reg_o >> 272; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "10";
            next_sm_specific_mac_address_b <= "10";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_12 =>
            -- -- In case of size 4
            -- reg_a = a0_0; reg_b = a2_0; reg_acc = reg_o; o2_0 = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "10";
            next_sm_specific_mac_address_o <= "10";
            next_sm_specific_mac_next_address_o <= "11";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_13 =>
            -- reg_a = a2_0; reg_b = a1_0; reg_acc = reg_o >> 272; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "10";
            next_sm_specific_mac_address_b <= "01";
            next_sm_specific_mac_address_o <= "11";
            next_sm_specific_mac_next_address_o <= "00";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_14 =>
            -- reg_a = a3_0; reg_b = a0_0; reg_acc = reg_o; o3_0 = reg_o; operation : 2*a*b + acc; Enable sign a; Increment o3_0 base address
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "11";
            next_sm_specific_mac_address_b <= "00";
            next_sm_specific_mac_address_o <= "11";
            next_sm_specific_mac_next_address_o <= "00";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '1';
        when square_direct_15 =>
            -- reg_a = a2_0; reg_b = a2_0; reg_acc = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "10";
            next_sm_specific_mac_address_b <= "10";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_16 =>
            -- reg_a = a3_0; reg_b = a1_0; reg_acc = reg_o; o4_0 = reg_o; Enable sign a; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "11";
            next_sm_specific_mac_address_b <= "01";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_17 =>
            -- reg_a = a3_0; reg_b = a2_0; reg_acc = reg_o >> 272; o5_0 = reg_o; Enable sign a; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "11";
            next_sm_specific_mac_address_b <= "10";
            next_sm_specific_mac_address_o <= "01";
            next_sm_specific_mac_next_address_o <= "10";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_direct_18 =>
            -- reg_a = a3_0; reg_b = a3_0; reg_acc = reg_o >> 272; o6_0 = reg_o; o7_0 = reg_o >> 272; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "11";
            next_sm_specific_mac_address_b <= "11";
            next_sm_specific_mac_address_o <= "10";
            next_sm_specific_mac_next_address_o <= "11";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_0 =>
            -- -- In case of size 1
            -- reg_a = a0_0; reg_b = b0_0; reg_acc = 0; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "00";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_1 =>
            -- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o0_0 = reg_y; operation : keep accumulator;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "11";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "00";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "10";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "11";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '1';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_2 =>
            -- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "00";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "01";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_3 =>
            -- reg_a = 0; reg_b = 0; reg_acc = reg_o >> 272; o0_0 = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "00";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "11";
            next_mac_clear_reg_b <= '1';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_5 =>
            -- -- In case of sizes 2, 3, 4
            -- reg_a = a0_0; reg_b = b0_0; reg_acc = 0; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "00";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_6 =>
            -- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o0_0 = reg_y; operation : keep accumulator;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "11";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "00";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "10";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "11";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '1';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_7 =>
            -- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "00";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "01";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_8 =>
            -- -- In case of size 2
            -- reg_a = a0_0; reg_b = b1_0; reg_acc = reg_o >> 272; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "01";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_9 =>
            -- reg_a = o0_0; reg_b = prime1; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "01";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_10 =>
            -- reg_a = a1_0; reg_b = b0_0; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "01";
            next_sm_specific_mac_address_b <= "00";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_11 =>
            -- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o1_0 = reg_y; operation : keep accumulator;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "11";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "00";
            next_sm_specific_mac_address_o <= "01";
            next_sm_specific_mac_next_address_o <= "10";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "10";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "11";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '1';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_12 =>
            -- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "00";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "01";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_13 =>
            -- reg_a = a1_0; reg_b = b1_0; reg_acc = reg_o >> 272; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "01";
            next_sm_specific_mac_address_b <= "01";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_14 =>
            -- reg_a = o1_0; reg_b = prime1; reg_acc = reg_o; o0_0 = reg_o; o1_0 = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "01";
            next_sm_specific_mac_address_b <= "01";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_16 =>
            -- -- In case of sizes 3, 4
            -- reg_a = a0_0; reg_b = b1_0; reg_acc = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "01";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_17 =>
            -- reg_a = o0_0; reg_b = prime1; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "01";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_18 =>
            -- reg_a = a1_0; reg_b = b0_0; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "01";
            next_sm_specific_mac_address_b <= "00";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_19 =>
            -- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o1_0 = reg_y; operation : keep accumulator;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "11";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "00";
            next_sm_specific_mac_address_o <= "01";
            next_sm_specific_mac_next_address_o <= "10";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "10";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "11";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '1';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_20 =>
            -- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "00";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "01";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_21 =>
            -- -- In case of size 3
            -- reg_a = a0_0; reg_b = b2_0; reg_acc = reg_o >> 272; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "10";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_22 =>
            -- reg_a = o0_0; reg_b = prime2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "10";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_23 =>
            -- reg_a = a1_0; reg_b = b1_0; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "01";
            next_sm_specific_mac_address_b <= "01";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_24 =>
            -- reg_a = o1_0; reg_b = prime1; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "01";
            next_sm_specific_mac_address_b <= "01";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_25 =>
            -- reg_a = a2_0; reg_b = b0_0; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "10";
            next_sm_specific_mac_address_b <= "00";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_26 =>
            -- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o2_0 = reg_y; operation : keep accumulator;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "11";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "00";
            next_sm_specific_mac_address_o <= "10";
            next_sm_specific_mac_next_address_o <= "11";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "10";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "11";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '1';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_27 =>
            -- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "00";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "01";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_28 =>
            -- reg_a = a1_0; reg_b = b2_0; reg_acc = reg_o >> 272; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "01";
            next_sm_specific_mac_address_b <= "10";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_29 =>
            -- reg_a = o1_0; reg_b = prime2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "01";
            next_sm_specific_mac_address_b <= "10";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_30 =>
            -- reg_a = a2_0; reg_b = b1_0; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "10";
            next_sm_specific_mac_address_b <= "01";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_31 =>
            -- reg_a = o2_0; reg_b = prime1; reg_acc = reg_o; o0_0 = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "10";
            next_sm_specific_mac_address_b <= "01";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_32 =>
            -- reg_a = a2_0; reg_b = b2_0; reg_acc = reg_o >> 272; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "10";
            next_sm_specific_mac_address_b <= "10";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_33 =>
            -- reg_a = o2_0; reg_b = prime2; reg_acc = reg_o; o1_0 = reg_o; o2_0 = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "10";
            next_sm_specific_mac_address_b <= "10";
            next_sm_specific_mac_address_o <= "01";
            next_sm_specific_mac_next_address_o <= "10";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_35 =>
            -- -- In case of size 4
            -- reg_a = a0_0; reg_b = b2_0; reg_acc = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "10";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_36 =>
            -- reg_a = o0_0; reg_b = prime2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "10";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_37 =>
            -- reg_a = a1_0; reg_b = b1_0; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "01";
            next_sm_specific_mac_address_b <= "01";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_38 =>
            -- reg_a = o1_0; reg_b = prime1; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "01";
            next_sm_specific_mac_address_b <= "01";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_39 =>
            -- reg_a = a2_0; reg_b = b0_0; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "10";
            next_sm_specific_mac_address_b <= "00";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_40 =>
            -- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o2_0 = reg_y; operation : keep accumulator;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "11";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "00";
            next_sm_specific_mac_address_o <= "10";
            next_sm_specific_mac_next_address_o <= "11";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "10";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "11";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '1';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_41 =>
            -- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "00";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "01";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_42 =>
            -- reg_a = a0_0; reg_b = b3_0; reg_acc = reg_o >> 272; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "11";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_43 =>
            -- reg_a = o0_0; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "11";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_44 =>
            -- reg_a = a1_0; reg_b = b2_0; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "01";
            next_sm_specific_mac_address_b <= "10";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_45 =>
            -- reg_a = o1_0; reg_b = prime2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "01";
            next_sm_specific_mac_address_b <= "10";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_46 =>
            -- reg_a = a2_0; reg_b = b1_0; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "10";
            next_sm_specific_mac_address_b <= "01";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_47 =>
            -- reg_a = o2_0; reg_b = prime1; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "10";
            next_sm_specific_mac_address_b <= "01";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_48 =>
            -- reg_a = a3_0; reg_b = b0_0; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "11";
            next_sm_specific_mac_address_b <= "00";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_49 =>
            -- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o3_0 = reg_y; operation : keep accumulator;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "11";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "00";
            next_sm_specific_mac_address_o <= "11";
            next_sm_specific_mac_next_address_o <= "00";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "10";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "11";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '1';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_50 =>
            -- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "00";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "01";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_51 =>
            -- reg_a = a1_0; reg_b = b3_0; reg_acc = reg_o >> 272; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "01";
            next_sm_specific_mac_address_b <= "11";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_52 =>
            -- reg_a = o1_0; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "01";
            next_sm_specific_mac_address_b <= "11";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_53 =>
            -- reg_a = a2_0; reg_b = b2_0; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "10";
            next_sm_specific_mac_address_b <= "10";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_54 =>
            -- reg_a = o2_0; reg_b = prime2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "10";
            next_sm_specific_mac_address_b <= "10";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_55 =>
            -- reg_a = a3_0; reg_b = b1_0; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "11";
            next_sm_specific_mac_address_b <= "01";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_56 =>
            -- reg_a = o3_0; reg_b = prime1; reg_acc = reg_o; o0_0 = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "11";
            next_sm_specific_mac_address_b <= "01";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_57 =>
            -- reg_a = a2_0; reg_b = b3_0; reg_acc = reg_o >> 272; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "10";
            next_sm_specific_mac_address_b <= "11";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_58 =>
            -- reg_a = o2_0; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "10";
            next_sm_specific_mac_address_b <= "11";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_59 =>
            -- reg_a = a3_0; reg_b = b2_0; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "11";
            next_sm_specific_mac_address_b <= "10";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_60 =>
            -- reg_a = o3_0; reg_b = prime2; reg_acc = reg_o; o1_0 = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "11";
            next_sm_specific_mac_address_b <= "10";
            next_sm_specific_mac_address_o <= "01";
            next_sm_specific_mac_next_address_o <= "10";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_61 =>
            -- reg_a = a3_0; reg_b = b3_0; reg_acc = reg_o >> 272; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "11";
            next_sm_specific_mac_address_b <= "11";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_62 =>
            -- reg_a = o3_0; reg_b = prime3; reg_acc = reg_o; o2_0 = reg_o; o3_0 = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "11";
            next_sm_specific_mac_address_b <= "11";
            next_sm_specific_mac_address_o <= "10";
            next_sm_specific_mac_next_address_o <= "11";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_0 =>
            -- -- In case of size 1
            -- reg_a = a0_0; reg_b = b0_0; reg_acc = 0; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "00";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_1 =>
            -- reg_a = 0; reg_b = 0; reg_acc = reg_o >> 272; o0_0 = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "00";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "11";
            next_mac_clear_reg_b <= '1';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_3 =>
            -- -- In case of sizes 2, 3, 4
            -- reg_a = a0_0; reg_b = b0_0; reg_acc = 0; o0_0 = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "00";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_4 =>
            -- -- In case of size 2
            -- reg_a = a0_0; reg_b = b1_0; reg_acc = reg_o >> 272; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "01";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_5 =>
            -- reg_a = o0_0; reg_b = primeSP1; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "01";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_6 =>
            -- reg_a = a1_0; reg_b = b0_0; reg_acc = reg_o; o1_0 = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "01";
            next_sm_specific_mac_address_b <= "00";
            next_sm_specific_mac_address_o <= "01";
            next_sm_specific_mac_next_address_o <= "10";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_7 =>
            -- reg_a = a1_0; reg_b = b1_0; reg_acc = reg_o >> 272; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "01";
            next_sm_specific_mac_address_b <= "01";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_8 =>
            -- reg_a = o1_0; reg_b = primeSP1; reg_acc = reg_o; o0_0 = reg_o; o1_0 = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "01";
            next_sm_specific_mac_address_b <= "01";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_10 =>
            -- -- In case of sizes 3, 4
            -- reg_a = a0_0; reg_b = b1_0; reg_acc = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "01";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_11 =>
            -- reg_a = o0_0; reg_b = primeSP1; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "01";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_12 =>
            -- reg_a = a1_0; reg_b = b0_0; reg_acc = reg_o; o1_0 = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "01";
            next_sm_specific_mac_address_b <= "00";
            next_sm_specific_mac_address_o <= "01";
            next_sm_specific_mac_next_address_o <= "10";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_13 =>
            -- -- In case of size 3
            -- reg_a = a0_0; reg_b = b2_0; reg_acc = reg_o >> 272; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "10";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_14 =>
            -- reg_a = o0_0; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "10";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_15 =>
            -- reg_a = a1_0; reg_b = b1_0; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "01";
            next_sm_specific_mac_address_b <= "01";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_16 =>
            -- reg_a = o1_0; reg_b = primeSP1; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "01";
            next_sm_specific_mac_address_b <= "01";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_17 =>
            -- reg_a = a2_0; reg_b = b0_0; reg_acc = reg_o; o2_0 = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "10";
            next_sm_specific_mac_address_b <= "00";
            next_sm_specific_mac_address_o <= "10";
            next_sm_specific_mac_next_address_o <= "11";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_18 =>
            -- reg_a = a1_0; reg_b = b2_0; reg_acc = reg_o >> 272; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "01";
            next_sm_specific_mac_address_b <= "10";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_19 =>
            -- reg_a = o1_0; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "01";
            next_sm_specific_mac_address_b <= "10";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_20 =>
            -- reg_a = a2_0; reg_b = b1_0; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "10";
            next_sm_specific_mac_address_b <= "01";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_21 =>
            -- reg_a = o2_0; reg_b = primeSP1; reg_acc = reg_o; o0_0 = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "10";
            next_sm_specific_mac_address_b <= "01";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_22 =>
            -- reg_a = a2_0; reg_b = b2_0; reg_acc = reg_o >> 272; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "10";
            next_sm_specific_mac_address_b <= "10";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_23 =>
            -- reg_a = o2_0; reg_b = primeSP2; reg_acc = reg_o; o1_0 = reg_o; o2_0 = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "10";
            next_sm_specific_mac_address_b <= "10";
            next_sm_specific_mac_address_o <= "01";
            next_sm_specific_mac_next_address_o <= "10";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_25 =>
            -- -- In case of size 4
            -- reg_a = a0_0; reg_b = b2_0; reg_acc = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "10";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_26 =>
            -- reg_a = o0_0; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "10";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_27 =>
            -- reg_a = a1_0; reg_b = b1_0; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "01";
            next_sm_specific_mac_address_b <= "01";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_28 =>
            -- reg_a = o1_0; reg_b = primeSP1; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "01";
            next_sm_specific_mac_address_b <= "01";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_29 =>
            -- reg_a = a2_0; reg_b = b0_0; reg_acc = reg_o; o2_0 = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "10";
            next_sm_specific_mac_address_b <= "00";
            next_sm_specific_mac_address_o <= "10";
            next_sm_specific_mac_next_address_o <= "11";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_30 =>
            -- reg_a = a0_0; reg_b = b3_0; reg_acc = reg_o >> 272; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "11";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_31 =>
            -- reg_a = o0_0; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "11";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_32 =>
            -- reg_a = a1_0; reg_b = b2_0; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "01";
            next_sm_specific_mac_address_b <= "10";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_33 =>
            -- reg_a = o1_0; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "01";
            next_sm_specific_mac_address_b <= "10";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_34 =>
            -- reg_a = a2_0; reg_b = b1_0; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "10";
            next_sm_specific_mac_address_b <= "01";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_35 =>
            -- reg_a = o2_0; reg_b = primeSP1; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "10";
            next_sm_specific_mac_address_b <= "01";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_36 =>
            -- reg_a = a3_0; reg_b = b0_0; reg_acc = reg_o; o3_0 = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "11";
            next_sm_specific_mac_address_b <= "00";
            next_sm_specific_mac_address_o <= "11";
            next_sm_specific_mac_next_address_o <= "00";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_37 =>
            -- reg_a = a1_0; reg_b = b3_0; reg_acc = reg_o >> 272; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "01";
            next_sm_specific_mac_address_b <= "11";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_38 =>
            -- reg_a = o1_0; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "01";
            next_sm_specific_mac_address_b <= "11";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_39 =>
            -- reg_a = a2_0; reg_b = b2_0; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "10";
            next_sm_specific_mac_address_b <= "10";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_40 =>
            -- reg_a = o2_0; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "10";
            next_sm_specific_mac_address_b <= "10";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_41 =>
            -- reg_a = a3_0; reg_b = b1_0; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "11";
            next_sm_specific_mac_address_b <= "01";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_42 =>
            -- reg_a = o3_0; reg_b = primeSP1; reg_acc = reg_o; o0_0 = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "11";
            next_sm_specific_mac_address_b <= "01";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_43 =>
            -- reg_a = a2_0; reg_b = b3_0; reg_acc = reg_o >> 272; Enable sign b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "10";
            next_sm_specific_mac_address_b <= "11";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_44 =>
            -- reg_a = o2_0; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "10";
            next_sm_specific_mac_address_b <= "11";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_45 =>
            -- reg_a = a3_0; reg_b = b2_0; reg_acc = reg_o; Enable sign a; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "11";
            next_sm_specific_mac_address_b <= "10";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_46 =>
            -- reg_a = o3_0; reg_b = primeSP2; reg_acc = reg_o; o1_0 = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "11";
            next_sm_specific_mac_address_b <= "10";
            next_sm_specific_mac_address_o <= "01";
            next_sm_specific_mac_next_address_o <= "10";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_47 =>
            -- reg_a = a3_0; reg_b = b3_0; reg_acc = reg_o >> 272; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "11";
            next_sm_specific_mac_address_b <= "11";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when multiplication_with_reduction_special_prime_48 =>
            -- reg_a = o3_0; reg_b = primeSP3; reg_acc = reg_o; o2_0 = reg_o; o3_0 = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "11";
            next_sm_specific_mac_address_b <= "11";
            next_sm_specific_mac_address_o <= "10";
            next_sm_specific_mac_next_address_o <= "11";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_0 =>
            -- -- In case of size 1
            -- reg_a = a0_0; reg_b = a0_0; reg_acc = 0; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "00";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_1 =>
            -- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o0_0 = reg_y; operation : keep accumulator;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "11";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "00";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "10";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "11";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '1';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_2 =>
            -- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "00";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "01";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_3 =>
            -- reg_a = 0; reg_b = 0; reg_acc = reg_o >> 272; o0_0 = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "00";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "11";
            next_mac_clear_reg_b <= '1';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_5 =>
            -- -- In case of 2, 3, 4
            -- reg_a = a0_0; reg_b = a0_0; reg_acc = 0; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "00";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_6 =>
            -- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o0_0 = reg_y; operation : keep accumulator;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "11";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "00";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "10";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "11";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '1';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_7 =>
            -- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "00";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "01";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_8 =>
            -- -- In case of size 2
            -- reg_a = a0_0; reg_b = a1_0; reg_acc = reg_o >> 272; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "01";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_9 =>
            -- reg_a = o0_0; reg_b = prime1; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "01";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_10 =>
            -- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o1_0 = reg_y; operation : keep accumulator;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "11";
            next_sm_specific_mac_address_a <= "01";
            next_sm_specific_mac_address_b <= "00";
            next_sm_specific_mac_address_o <= "01";
            next_sm_specific_mac_next_address_o <= "10";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "10";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "11";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '1';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_11 =>
            -- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "01";
            next_sm_specific_mac_address_b <= "00";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "01";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_12 =>
            -- reg_a = a1_0; reg_b = a1_0; reg_acc = reg_o >> 272; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "01";
            next_sm_specific_mac_address_b <= "01";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_13 =>
            -- reg_a = o1_0; reg_b = prime1; reg_acc = reg_o; o0_0 = reg_o; o1_0 = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "01";
            next_sm_specific_mac_address_b <= "01";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_15 =>
            -- -- In case of size 3, 4
            -- reg_a = a0_0; reg_b = a1_0; reg_acc = reg_o >> 272; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "01";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_16 =>
            -- reg_a = o0_0; reg_b = prime1; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "01";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_17 =>
            -- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o1_0 = reg_y; operation : keep accumulator;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "11";
            next_sm_specific_mac_address_a <= "01";
            next_sm_specific_mac_address_b <= "00";
            next_sm_specific_mac_address_o <= "01";
            next_sm_specific_mac_next_address_o <= "10";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "10";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "11";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '1';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_18 =>
            -- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "01";
            next_sm_specific_mac_address_b <= "00";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "01";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_19 =>
            -- -- In case of size 3
            -- reg_a = a0_0; reg_b = a2_0; reg_acc = reg_o >> 272; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "10";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_20 =>
            -- reg_a = o0_0; reg_b = prime2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "10";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_21 =>
            -- reg_a = a1_0; reg_b = a1_0; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "01";
            next_sm_specific_mac_address_b <= "01";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_22 =>
            -- reg_a = o1_0; reg_b = prime1; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "01";
            next_sm_specific_mac_address_b <= "01";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_23 =>
            -- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o2_0 = reg_y; operation : keep accumulator;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "11";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "00";
            next_sm_specific_mac_address_o <= "10";
            next_sm_specific_mac_next_address_o <= "11";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "10";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "11";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '1';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_24 =>
            -- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "00";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "01";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_25 =>
            -- reg_a = a1_0; reg_b = a2_0; reg_acc = reg_o >> 272; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "01";
            next_sm_specific_mac_address_b <= "10";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_26 =>
            -- reg_a = o1_0; reg_b = prime2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "01";
            next_sm_specific_mac_address_b <= "10";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_27 =>
            -- reg_a = o2_0; reg_b = prime1; reg_acc = reg_o; o0_0 = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "10";
            next_sm_specific_mac_address_b <= "01";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_28 =>
            -- reg_a = a2_0; reg_b = a2_0; reg_acc = reg_o >> 272; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "10";
            next_sm_specific_mac_address_b <= "10";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_29 =>
            -- reg_a = o2_0; reg_b = prime2; reg_acc = reg_o; o1_0 = reg_o; o2_0 = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "10";
            next_sm_specific_mac_address_b <= "10";
            next_sm_specific_mac_address_o <= "01";
            next_sm_specific_mac_next_address_o <= "10";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_31 =>
            -- -- In case of size 4
            -- reg_a = a0_0; reg_b = a2_0; reg_acc = reg_o >> 272; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "10";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_32 =>
            -- reg_a = o0_0; reg_b = prime2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "10";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_33 =>
            -- reg_a = a1_0; reg_b = a1_0; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "01";
            next_sm_specific_mac_address_b <= "01";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_34 =>
            -- reg_a = o1_0; reg_b = prime1; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "01";
            next_sm_specific_mac_address_b <= "01";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_35 =>
            -- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o2_0 = reg_y; operation : keep accumulator;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "11";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "00";
            next_sm_specific_mac_address_o <= "10";
            next_sm_specific_mac_next_address_o <= "11";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "10";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "11";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '1';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_36 =>
            -- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "00";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "01";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_37 =>
            -- reg_a = a0_0; reg_b = a3_0; reg_acc = reg_o >> 272; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "11";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_38 =>
            -- reg_a = o0_0; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "11";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_39 =>
            -- reg_a = a1_0; reg_b = a2_0; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "01";
            next_sm_specific_mac_address_b <= "10";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_40 =>
            -- reg_a = o1_0; reg_b = prime2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "01";
            next_sm_specific_mac_address_b <= "10";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_41 =>
            -- reg_a = o2_0; reg_b = prime1; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "10";
            next_sm_specific_mac_address_b <= "01";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_42 =>
            -- reg_a = reg_o; reg_b = prime_line_0; reg_acc = reg_o; o3_0 = reg_y; operation : keep accumulator;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "11";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "00";
            next_sm_specific_mac_address_o <= "11";
            next_sm_specific_mac_next_address_o <= "00";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "10";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "11";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '1';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_43 =>
            -- reg_a = reg_y; reg_b = prime0; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "00";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "01";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_44 =>
            -- reg_a = a1_0; reg_b = a3_0; reg_acc = reg_o >> 272; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "01";
            next_sm_specific_mac_address_b <= "11";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_45 =>
            -- reg_a = o1_0; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "01";
            next_sm_specific_mac_address_b <= "11";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_46 =>
            -- reg_a = a2_0; reg_b = a2_0; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "10";
            next_sm_specific_mac_address_b <= "10";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_47 =>
            -- reg_a = o2_0; reg_b = prime2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "10";
            next_sm_specific_mac_address_b <= "10";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_48 =>
            -- reg_a = o3_0; reg_b = prime1; reg_acc = reg_o; o0_0 = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "11";
            next_sm_specific_mac_address_b <= "01";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_49 =>
            -- reg_a = a2_0; reg_b = a3_0; reg_acc = reg_o >> 272; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "10";
            next_sm_specific_mac_address_b <= "11";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_50 =>
            -- reg_a = o2_0; reg_b = prime3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "10";
            next_sm_specific_mac_address_b <= "11";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_51 =>
            -- reg_a = o3_0; reg_b = prime2; reg_acc = reg_o; o1_0 = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "11";
            next_sm_specific_mac_address_b <= "10";
            next_sm_specific_mac_address_o <= "01";
            next_sm_specific_mac_next_address_o <= "10";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_52 =>
            -- reg_a = a3_0; reg_b = a3_0; reg_acc = reg_o >> 272; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "11";
            next_sm_specific_mac_address_b <= "11";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_53 =>
            -- reg_a = o3_0; reg_b = prime3; reg_acc = reg_o; o2_0 = reg_o; o3_0 = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "11";
            next_sm_specific_mac_address_b <= "11";
            next_sm_specific_mac_address_o <= "10";
            next_sm_specific_mac_next_address_o <= "11";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_0 =>
            -- -- In case of size 1
            -- reg_a = a0_0; reg_b = a0_0; reg_acc = 0; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "00";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_1 =>
            -- reg_a = 0; reg_b = 0; reg_acc = reg_o >> 272; o0_0 = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "00";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "11";
            next_mac_clear_reg_b <= '1';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_3 =>
            -- -- In case of size 2, 3, 4
            -- reg_a = a0_0; reg_b = a0_0; reg_acc = 0; o0_0 = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "00";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_4 =>
            -- -- In case of size 2
            -- reg_a = a0_0; reg_b = a1_0; reg_acc = reg_o >> 272; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "01";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_5 =>
            -- reg_a = o0_0; reg_b = primeSP1; reg_acc = reg_o; o1_0 = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "01";
            next_sm_specific_mac_address_o <= "01";
            next_sm_specific_mac_next_address_o <= "10";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_6 =>
            -- reg_a = a1_0; reg_b = a1_0; reg_acc = reg_o >> 272; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "01";
            next_sm_specific_mac_address_b <= "01";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_7 =>
            -- reg_a = o1_0; reg_b = primeSP1; reg_acc = reg_o; o0_0 = reg_o; o1_0 = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "01";
            next_sm_specific_mac_address_b <= "01";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_9 =>
            -- -- In case of size 3, 4
            -- reg_a = a0_0; reg_b = a1_0; reg_acc = reg_o >> 272; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "01";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_10 =>
            -- reg_a = o0_0; reg_b = primeSP1; reg_acc = reg_o; o1_0 = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "01";
            next_sm_specific_mac_address_o <= "01";
            next_sm_specific_mac_next_address_o <= "10";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_11 =>
            -- -- In case of size 3
            -- reg_a = a0_0; reg_b = a2_0; reg_acc = reg_o >> 272; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "10";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_12 =>
            -- reg_a = o0_0; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "10";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_13 =>
            -- reg_a = a1_0; reg_b = a1_0; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "01";
            next_sm_specific_mac_address_b <= "01";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_14 =>
            -- reg_a = o1_0; reg_b = primeSP1; reg_acc = reg_o; o2_0 = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "01";
            next_sm_specific_mac_address_b <= "01";
            next_sm_specific_mac_address_o <= "10";
            next_sm_specific_mac_next_address_o <= "11";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_15 =>
            -- reg_a = a1_0; reg_b = a2_0; reg_acc = reg_o >> 272; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "01";
            next_sm_specific_mac_address_b <= "10";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_16 =>
            -- reg_a = o1_0; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "01";
            next_sm_specific_mac_address_b <= "10";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_17 =>
            -- reg_a = o2_0; reg_b = primeSP1; reg_acc = reg_o; o0_0 = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "10";
            next_sm_specific_mac_address_b <= "01";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_18 =>
            -- reg_a = a2_0; reg_b = a2_0; reg_acc = reg_o >> 272; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "10";
            next_sm_specific_mac_address_b <= "10";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_19 =>
            -- reg_a = o2_0; reg_b = primeSP2; reg_acc = reg_o; o1_0 = reg_o; o2_0 = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "10";
            next_sm_specific_mac_address_b <= "10";
            next_sm_specific_mac_address_o <= "01";
            next_sm_specific_mac_next_address_o <= "10";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_21 =>
            -- -- In case of size 4
            -- reg_a = a0_0; reg_b = a2_0; reg_acc = reg_o >> 272; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "10";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_22 =>
            -- reg_a = o0_0; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "10";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_23 =>
            -- reg_a = a1_0; reg_b = a1_0; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "01";
            next_sm_specific_mac_address_b <= "01";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_24 =>
            -- reg_a = o1_0; reg_b = primeSP1; reg_acc = reg_o; o2_0 = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "01";
            next_sm_specific_mac_address_b <= "01";
            next_sm_specific_mac_address_o <= "10";
            next_sm_specific_mac_next_address_o <= "11";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_25 =>
            -- reg_a = a0_0; reg_b = a3_0; reg_acc = reg_o >> 272; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "11";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_26 =>
            -- reg_a = o0_0; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "11";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_27 =>
            -- reg_a = a1_0; reg_b = a2_0; reg_acc = reg_o; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "01";
            next_sm_specific_mac_address_b <= "10";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_28 =>
            -- reg_a = o1_0; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "01";
            next_sm_specific_mac_address_b <= "10";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_29 =>
            -- reg_a = o2_0; reg_b = primeSP1; reg_acc = reg_o; o3_0 = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "10";
            next_sm_specific_mac_address_b <= "01";
            next_sm_specific_mac_address_o <= "11";
            next_sm_specific_mac_next_address_o <= "00";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_30 =>
            -- reg_a = a1_0; reg_b = a3_0; reg_acc = reg_o >> 272; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "01";
            next_sm_specific_mac_address_b <= "11";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_31 =>
            -- reg_a = o1_0; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "01";
            next_sm_specific_mac_address_b <= "11";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_32 =>
            -- reg_a = a2_0; reg_b = a2_0; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "10";
            next_sm_specific_mac_address_b <= "10";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_33 =>
            -- reg_a = o2_0; reg_b = primeSP2; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "10";
            next_sm_specific_mac_address_b <= "10";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_34 =>
            -- reg_a = o3_0; reg_b = primeSP1; reg_acc = reg_o; o0_0 = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "11";
            next_sm_specific_mac_address_b <= "01";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_35 =>
            -- reg_a = a2_0; reg_b = a3_0; reg_acc = reg_o >> 272; Enable sign b; operation : 2*a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "10";
            next_sm_specific_mac_address_b <= "11";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '1';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_36 =>
            -- reg_a = o2_0; reg_b = primeSP3; reg_acc = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "10";
            next_sm_specific_mac_address_b <= "11";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_37 =>
            -- reg_a = o3_0; reg_b = primeSP2; reg_acc = reg_o; o1_0 = reg_o; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "11";
            next_sm_specific_mac_address_b <= "10";
            next_sm_specific_mac_address_o <= "01";
            next_sm_specific_mac_next_address_o <= "10";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_38 =>
            -- reg_a = a3_0; reg_b = a3_0; reg_acc = reg_o >> 272; Enable sign a,b; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "11";
            next_sm_specific_mac_address_b <= "11";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when square_with_reduction_special_prime_39 =>
            -- reg_a = o3_0; reg_b = primeSP3; reg_acc = reg_o; o2_0 = reg_o; o3_0 = reg_o >> 272; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "11";
            next_sm_specific_mac_address_b <= "11";
            next_sm_specific_mac_address_o <= "10";
            next_sm_specific_mac_next_address_o <= "11";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '1';
            next_mac_memory_only_write_mode <= '1';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_direct_0 =>
            -- -- In case of size 1
            -- reg_a = a0_0; reg_b = b0_0; reg_acc = 0; o0_0 = reg_o; Enable sign a,b; operation : b +/- a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "00";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '1';
            next_sm_mac_operation_mode(1) <= '0';
            next_sm_mac_operation_mode(0) <= '0';
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_direct_2 =>
            -- -- In case of size 2, 3, 4
            -- reg_a = a0_0; reg_b = b0_0; reg_acc = 0; o0_0 = reg_o; operation : b +/- a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "00";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '1';
            next_sm_mac_operation_mode(1) <= '0';
            next_sm_mac_operation_mode(0) <= '0';
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_direct_3 =>
            -- -- In case of size 2
            -- reg_a = a1_0; reg_b = b1_0; reg_acc = reg_o >> 272; o1_0 = reg_o; Enable sign a,b; operation : b +/- a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "01";
            next_sm_specific_mac_address_b <= "01";
            next_sm_specific_mac_address_o <= "01";
            next_sm_specific_mac_next_address_o <= "10";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '1';
            next_sm_mac_operation_mode(1) <= '0';
            next_sm_mac_operation_mode(0) <= '0';
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_direct_5 =>
            -- -- In case of size 3, 4
            -- reg_a = a1_0; reg_b = b1_0; reg_acc = reg_o >> 272; o1_0 = reg_o; operation : b +/- a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "01";
            next_sm_specific_mac_address_b <= "01";
            next_sm_specific_mac_address_o <= "01";
            next_sm_specific_mac_next_address_o <= "10";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '1';
            next_sm_mac_operation_mode(1) <= '0';
            next_sm_mac_operation_mode(0) <= '0';
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_direct_6 =>
            -- -- In case of size 3
            -- reg_a = a2_0; reg_b = b2_0; reg_acc = reg_o >> 272; o2_0 = reg_o; Enable sign a,b; operation : b +/- a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "10";
            next_sm_specific_mac_address_b <= "10";
            next_sm_specific_mac_address_o <= "10";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '1';
            next_sm_mac_operation_mode(1) <= '0';
            next_sm_mac_operation_mode(0) <= '0';
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_direct_8 =>
            -- -- In case of size 4
            -- reg_a = a2_0; reg_b = b2_0; reg_acc = reg_o >> 272; o2_0 = reg_o; operation : b +/- a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "10";
            next_sm_specific_mac_address_b <= "10";
            next_sm_specific_mac_address_o <= "10";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '1';
            next_sm_mac_operation_mode(1) <= '0';
            next_sm_mac_operation_mode(0) <= '0';
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when addition_subtraction_direct_9 =>
            -- reg_a = a3_0; reg_b = b3_0; reg_acc = reg_o >> 272; o3_0 = reg_o; Enable sign a,b; operation : b +/- a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "11";
            next_sm_specific_mac_address_b <= "11";
            next_sm_specific_mac_address_o <= "11";
            next_sm_specific_mac_next_address_o <= "00";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '1';
            next_sm_mac_operation_mode(1) <= '0';
            next_sm_mac_operation_mode(0) <= '0';
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_0 =>
            -- reg_a = a0_0; reg_b = 0; reg_acc = 0; Enable sign a,b; operation : b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "00";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '1';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_1 =>
            -- reg_a = 0; reg_b = prime_0; reg_acc = reg_o; reg_s = reg_o_positive; Enable sign a,b; operation : -s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "00";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "11";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '1';
            next_mac_sel_reg_s_reg_o_sign <= '1';
            next_mac_reg_s_reg_o_positive <= '1';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_2 =>
            -- reg_a = 0; reg_b = prime_0; reg_acc = reg_o; reg_s = reg_o_negative; Enable sign a,b; operation : s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "00";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "11";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '1';
            next_mac_sel_reg_s_reg_o_sign <= '1';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_3 =>
            -- reg_a = 0; reg_b = prime_0; reg_acc = reg_o; o0_0 = reg_o; reg_s = reg_o_negative; Enable sign a,b; operation : s*b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "00";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "11";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '1';
            next_mac_sel_reg_s_reg_o_sign <= '1';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_5 =>
            -- reg_a = a1_0; reg_b = 0; reg_acc = 0; Enable sign a,b; operation : b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "01";
            next_sm_specific_mac_address_b <= "00";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '1';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_6 =>
            -- reg_a = a0_0; reg_b = prime_0; reg_acc = 0; o0_0 = reg_o; reg_s = reg_o_positive; operation : -s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "00";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '1';
            next_mac_sel_reg_s_reg_o_sign <= '1';
            next_mac_reg_s_reg_o_positive <= '1';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_7 =>
            -- reg_a = a1_0; reg_b = prime_1; reg_acc = reg_o >> 272; o1_0 = reg_o; Enable sign a,b; operation : -s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "01";
            next_sm_specific_mac_address_b <= "01";
            next_sm_specific_mac_address_o <= "01";
            next_sm_specific_mac_next_address_o <= "10";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_8 =>
            -- reg_a = o0_0; reg_b = prime_0; reg_acc = 0; o0_0 = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "00";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '1';
            next_mac_sel_reg_s_reg_o_sign <= '1';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_9 =>
            -- reg_a = o1_0; reg_b = prime_1; reg_acc = reg_o >> 272; o1_0 = reg_o; Enable sign a,b operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "01";
            next_sm_specific_mac_address_b <= "01";
            next_sm_specific_mac_address_o <= "01";
            next_sm_specific_mac_next_address_o <= "10";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_10 =>
            -- reg_a = o0_0; reg_b = prime_0; reg_acc = 0; o0_0 = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "00";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '1';
            next_mac_sel_reg_s_reg_o_sign <= '1';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_11 =>
            -- reg_a = o1_0; reg_b = prime_1; reg_acc = reg_o >> 272; o1_0 = reg_o; Enable sign a,b operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "01";
            next_sm_specific_mac_address_b <= "01";
            next_sm_specific_mac_address_o <= "01";
            next_sm_specific_mac_next_address_o <= "10";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_13 =>
            -- reg_a = a2_0; reg_b = 0; reg_acc = 0; Enable sign a,b; operation : b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "10";
            next_sm_specific_mac_address_b <= "10";
            next_sm_specific_mac_address_o <= "10";
            next_sm_specific_mac_next_address_o <= "11";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '1';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_14 =>
            -- reg_a = a0_0; reg_b = prime_0; reg_acc = 0; o0_0 = reg_o; reg_s = reg_o_positive; operation : -s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "00";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '1';
            next_mac_sel_reg_s_reg_o_sign <= '1';
            next_mac_reg_s_reg_o_positive <= '1';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_15 =>
            -- reg_a = a1_0; reg_b = prime_1; reg_acc = reg_o >> 272; o1_0 = reg_o; operation : -s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "01";
            next_sm_specific_mac_address_b <= "01";
            next_sm_specific_mac_address_o <= "01";
            next_sm_specific_mac_next_address_o <= "10";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_16 =>
            -- reg_a = a2_0; reg_b = prime_2; reg_acc = reg_o >> 272; o2_0 = reg_o; Enable sign a,b; operation : -s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "10";
            next_sm_specific_mac_address_b <= "10";
            next_sm_specific_mac_address_o <= "10";
            next_sm_specific_mac_next_address_o <= "11";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_17 =>
            -- reg_a = o0_0; reg_b = prime_0; reg_acc = 0; o0_0 = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "00";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '1';
            next_mac_sel_reg_s_reg_o_sign <= '1';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_18 =>
            -- reg_a = o1_0; reg_b = prime_1; reg_acc = reg_o >> 272; o1_0 = reg_o; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "01";
            next_sm_specific_mac_address_b <= "01";
            next_sm_specific_mac_address_o <= "01";
            next_sm_specific_mac_next_address_o <= "10";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_19 =>
            -- reg_a = o2_0; reg_b = prime_2; reg_acc = reg_o >> 272; o2_0 = reg_o; Enable sign a,b operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "10";
            next_sm_specific_mac_address_b <= "10";
            next_sm_specific_mac_address_o <= "10";
            next_sm_specific_mac_next_address_o <= "11";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_20 =>
            -- reg_a = o0_0; reg_b = prime_0; reg_acc = 0; o0_0 = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "00";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '1';
            next_mac_sel_reg_s_reg_o_sign <= '1';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_21 =>
            -- reg_a = o1_0; reg_b = prime_1; reg_acc = reg_o >> 272; o1_0 = reg_o; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "01";
            next_sm_specific_mac_address_b <= "01";
            next_sm_specific_mac_address_o <= "01";
            next_sm_specific_mac_next_address_o <= "10";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_22 =>
            -- reg_a = o2_0; reg_b = prime_2; reg_acc = reg_o >> 272; o2_0 = reg_o; Enable sign a,b operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "10";
            next_sm_specific_mac_address_b <= "10";
            next_sm_specific_mac_address_o <= "10";
            next_sm_specific_mac_next_address_o <= "11";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_24 =>
            -- reg_a = a3_0; reg_b = 0; reg_acc = 0; Enable sign a,b; operation : b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "11";
            next_sm_specific_mac_address_b <= "11";
            next_sm_specific_mac_address_o <= "11";
            next_sm_specific_mac_next_address_o <= "00";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '1';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_25 =>
            -- reg_a = a0_0; reg_b = prime_0; reg_acc = 0; o0_0 = reg_o; reg_s = reg_o_positive; operation : -s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "00";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '1';
            next_mac_sel_reg_s_reg_o_sign <= '1';
            next_mac_reg_s_reg_o_positive <= '1';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_26 =>
            -- reg_a = a1_0; reg_b = prime_1; reg_acc = reg_o >> 272; o1_0 = reg_o; operation : -s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "01";
            next_sm_specific_mac_address_b <= "01";
            next_sm_specific_mac_address_o <= "01";
            next_sm_specific_mac_next_address_o <= "10";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_27 =>
            -- reg_a = a2_0; reg_b = prime_2; reg_acc = reg_o >> 272; o2_0 = reg_o; operation : -s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "10";
            next_sm_specific_mac_address_b <= "10";
            next_sm_specific_mac_address_o <= "10";
            next_sm_specific_mac_next_address_o <= "11";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_28 =>
            -- reg_a = a3_0; reg_b = prime_3; reg_acc = reg_o >> 272; o3_0 = reg_o; Enable sign a,b; operation : -s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "11";
            next_sm_specific_mac_address_b <= "11";
            next_sm_specific_mac_address_o <= "11";
            next_sm_specific_mac_next_address_o <= "00";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "00";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '1';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_29 =>
            -- reg_a = o0_0; reg_b = prime_0; reg_acc = 0; o0_0 = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "00";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '1';
            next_mac_sel_reg_s_reg_o_sign <= '1';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_30 =>
            -- reg_a = o1_0; reg_b = prime_1; reg_acc = reg_o >> 272; o1_0 = reg_o; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "01";
            next_sm_specific_mac_address_b <= "01";
            next_sm_specific_mac_address_o <= "01";
            next_sm_specific_mac_next_address_o <= "10";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_31 =>
            -- reg_a = o2_0; reg_b = prime_2; reg_acc = reg_o >> 272; o2_0 = reg_o; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "10";
            next_sm_specific_mac_address_b <= "10";
            next_sm_specific_mac_address_o <= "10";
            next_sm_specific_mac_next_address_o <= "11";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_32 =>
            -- reg_a = o3_0; reg_b = prime_3; reg_acc = reg_o >> 272; o3_0 = reg_o; Enable sign a,b; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "11";
            next_sm_specific_mac_address_b <= "11";
            next_sm_specific_mac_address_o <= "11";
            next_sm_specific_mac_next_address_o <= "00";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_33 =>
            -- reg_a = o0_0; reg_b = prime_0; reg_acc = 0; o0_0 = reg_o; reg_s = reg_o_negative; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "00";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '1';
            next_mac_sel_reg_s_reg_o_sign <= '1';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_34 =>
            -- reg_a = o1_0; reg_b = prime_1; reg_acc = reg_o >> 272; o1_0 = reg_o; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "01";
            next_sm_specific_mac_address_b <= "01";
            next_sm_specific_mac_address_o <= "01";
            next_sm_specific_mac_next_address_o <= "10";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_35 =>
            -- reg_a = o2_0; reg_b = prime_2; reg_acc = reg_o >> 272; o2_0 = reg_o; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "10";
            next_sm_specific_mac_address_b <= "10";
            next_sm_specific_mac_address_o <= "10";
            next_sm_specific_mac_next_address_o <= "11";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when iterative_modular_reduction_36 =>
            -- reg_a = o3_0; reg_b = prime_3; reg_acc = reg_o >> 272; o3_0 = reg_o; Enable sign a,b; operation : s*b + a + acc
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '1';
            next_sel_address_b_prime <= "10";
            next_sm_specific_mac_address_a <= "11";
            next_sm_specific_mac_address_b <= "11";
            next_sm_specific_mac_address_o <= "11";
            next_sm_specific_mac_next_address_o <= "00";
            next_mac_enable_signed_a <= '1';
            next_mac_enable_signed_b <= '1';
            next_mac_sel_load_reg_a <= "00";
            next_mac_clear_reg_b <= '0';
            next_mac_clear_reg_acc <= '0';
            next_mac_sel_shift_reg_o <= '1';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '1';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '1';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when nop_4_stages =>
        -- reg_a = 0; reg_b = 0; reg_acc = 0; operation : b + a + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "10";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "00";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "11";
            next_mac_clear_reg_b <= '1';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "01";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
        when nop_8_stages =>
        -- reg_a = 0; reg_b = 0; reg_acc = 0; operation : a*b + acc;
            next_sm_free_flag <= '0';
            next_sm_rotation_size <= "11";
            next_sm_circular_shift_enable <= '1';
            next_sel_address_a <= '0';
            next_sel_address_b_prime <= "00";
            next_sm_specific_mac_address_a <= "00";
            next_sm_specific_mac_address_b <= "00";
            next_sm_specific_mac_address_o <= "00";
            next_sm_specific_mac_next_address_o <= "01";
            next_mac_enable_signed_a <= '0';
            next_mac_enable_signed_b <= '0';
            next_mac_sel_load_reg_a <= "11";
            next_mac_clear_reg_b <= '1';
            next_mac_clear_reg_acc <= '1';
            next_mac_sel_shift_reg_o <= '0';
            next_mac_enable_update_reg_s <= '0';
            next_mac_sel_reg_s_reg_o_sign <= '0';
            next_mac_reg_s_reg_o_positive <= '0';
            next_sm_sign_a_mode <= '0';
            next_sm_mac_operation_mode <= "10";
            next_mac_enable_reg_s_mask <= '0';
            next_mac_subtraction_reg_a_b <= '0';
            next_mac_sel_multiply_two_a_b <= '0';
            next_mac_sel_reg_y_output <= '0';
            next_sm_mac_write_enable_output <= '0';
            next_mac_memory_double_mode <= '0';
            next_mac_memory_only_write_mode <= '0';
            next_base_address_generator_o_increment_previous_address <= '0';
--        when others => 
--            next_sm_free_flag <= '0';
--            next_sm_rotation_size <= "11";
--            next_sm_circular_shift_enable <= '0';
--            next_sel_address_a <= '0';
--            next_sel_address_b_prime <= "00";
--            next_sm_specific_mac_address_a <= "00";
--            next_sm_specific_mac_address_b <= "00";
--            next_sm_specific_mac_address_o <= "00";
--            next_sm_specific_mac_next_address_o <= "01";
--            next_mac_enable_signed_a <= '0';
--            next_mac_enable_signed_b <= '0';
--            next_mac_sel_load_reg_a <= "11";
--            next_mac_clear_reg_b <= '1';
--            next_mac_clear_reg_acc <= '1';
--            next_mac_sel_shift_reg_o <= '0';
--            next_mac_enable_update_reg_s <= '0';
--            next_mac_sel_reg_s_reg_o_sign <= '0';
--            next_mac_reg_s_reg_o_positive <= '0';
--            next_sm_sign_a_mode <= '0';
--            next_sm_mac_operation_mode <= "10";
--            next_mac_enable_reg_s_mask <= '0';
--            next_mac_subtraction_reg_a_b <= '0';
--            next_mac_sel_multiply_two_a_b <= '0';
--            next_mac_sel_reg_y_output <= '0';
--            next_sm_mac_write_enable_output <= '0';
--            next_mac_memory_double_mode <= '0';
--            next_mac_memory_only_write_mode <= '0';
--            next_base_address_generator_o_increment_previous_address <= '0';
    end case;
end process;

update_state : process(actual_state, instruction_values_valid, instruction_type, prime_line_equal_one, operands_size, penultimate_operation)
begin
case (actual_state) is
        when reset =>
            next_state <= decode_instruction;
        when decode_instruction =>
            next_state <= decode_instruction;
            if(instruction_values_valid = '1') then
                if(instruction_type = "0000") then
                    if(operands_size = "00") then
                        next_state <= multiplication_direct_0;
                    else
                        next_state <= multiplication_direct_2;
                    end if;
                elsif(instruction_type = "0001") then
                    if(operands_size = "00") then
                        next_state <= square_direct_0;
                    else
                        next_state <= square_direct_2;
                    end if;
                elsif(instruction_type = "0010") then
                    if(prime_line_equal_one = '1') then
                        if(operands_size = "00") then
                            next_state <= multiplication_with_reduction_special_prime_0;
                        else
                            next_state <= multiplication_with_reduction_special_prime_3;
                        end if;
                    else
                        if(operands_size = "00") then
                            next_state <= multiplication_with_reduction_0;
                        else
                            next_state <= multiplication_with_reduction_5;
                        end if;
                    end if;
                elsif(instruction_type = "0011") then
                    if(prime_line_equal_one = '1') then
                        if(operands_size = "00") then
                            next_state <= square_with_reduction_special_prime_0;
                        else
                            next_state <= square_with_reduction_special_prime_3;
                        end if;
                    else
                        if(operands_size = "00") then
                            next_state <= square_with_reduction_0;
                        else
                            next_state <= square_with_reduction_5;
                        end if;
                    end if;
                elsif(instruction_type = "0100") then
                    if(operands_size = "00") then
                        next_state <= addition_subtraction_direct_0;
                    else
                        next_state <= addition_subtraction_direct_2;
                    end if;
                elsif(instruction_type = "0101") then
                    if(operands_size = "00") then
                        next_state <= iterative_modular_reduction_0;
                    elsif(operands_size = "01") then
                        next_state <= iterative_modular_reduction_5;
                    elsif(operands_size = "10") then
                        next_state <= iterative_modular_reduction_13;
                    else
                        next_state <= iterative_modular_reduction_24;
                    end if;
                end if;
            end if;
        when multiplication_direct_0 =>
            next_state <= multiplication_direct_0;
            if(penultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when multiplication_direct_2 =>
            next_state <= multiplication_direct_2;
            if(penultimate_operation = '1') then
                if(operands_size = "01") then
                    next_state <= multiplication_direct_3;
                else
                    next_state <= multiplication_direct_7;
                end if;
            end if;
        when multiplication_direct_3 =>
            next_state <= multiplication_direct_3;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_4;
            end if;
        when multiplication_direct_4 =>
            next_state <= multiplication_direct_4;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_5;
            end if;
        when multiplication_direct_5 =>
            next_state <= multiplication_direct_5;
            if(penultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when multiplication_direct_7 =>
            next_state <= multiplication_direct_7;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_8;
            end if;
        when multiplication_direct_8 =>
            next_state <= multiplication_direct_8;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_9;
            end if;
        when multiplication_direct_9 =>
            next_state <= multiplication_direct_9;
            if(penultimate_operation = '1') then
                if(operands_size = "10") then
                    next_state <= multiplication_direct_10;
                else
                    next_state <= multiplication_direct_16;
                end if;
            end if;
        when multiplication_direct_10 =>
            next_state <= multiplication_direct_10;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_11;
            end if;
        when multiplication_direct_11 =>
            next_state <= multiplication_direct_11;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_12;
            end if;
        when multiplication_direct_12 =>
            next_state <= multiplication_direct_12;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_13;
            end if;
        when multiplication_direct_13 =>
            next_state <= multiplication_direct_13;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_14;
            end if;
        when multiplication_direct_14 =>
            next_state <= multiplication_direct_14;
            if(penultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when multiplication_direct_16 =>
            next_state <= multiplication_direct_16;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_17;
            end if;
        when multiplication_direct_17 =>
            next_state <= multiplication_direct_17;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_18;
            end if;
        when multiplication_direct_18 =>
            next_state <= multiplication_direct_18;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_19;
            end if;
        when multiplication_direct_19 =>
            next_state <= multiplication_direct_19;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_20;
            end if;
        when multiplication_direct_20 =>
            next_state <= multiplication_direct_20;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_21;
            end if;
        when multiplication_direct_21 =>
            next_state <= multiplication_direct_21;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_22;
            end if;
        when multiplication_direct_22 =>
            next_state <= multiplication_direct_22;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_23;
            end if;
        when multiplication_direct_23 =>
            next_state <= multiplication_direct_23;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_24;
            end if;
        when multiplication_direct_24 =>
            next_state <= multiplication_direct_24;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_25;
            end if;
        when multiplication_direct_25 =>
            next_state <= multiplication_direct_25;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_26;
            end if;
        when multiplication_direct_26 =>
            next_state <= multiplication_direct_26;
            if(penultimate_operation = '1') then
                next_state <= multiplication_direct_27;
            end if;
        when multiplication_direct_27 =>
            next_state <= multiplication_direct_27;
            if(penultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when square_direct_0 => 
            next_state <= square_direct_0;
            if(penultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when square_direct_2 => 
            next_state <= square_direct_2;
            if(penultimate_operation = '1') then
                if(operands_size = "01") then
                    next_state <= square_direct_3;
                else
                    next_state <= square_direct_6;
                end if;
            end if;
        when square_direct_3 => 
            next_state <= square_direct_3;
            if(penultimate_operation = '1') then
                next_state <= square_direct_4;
            end if;
        when square_direct_4 => 
            next_state <= square_direct_4;
            if(penultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when square_direct_6 => 
            next_state <= square_direct_6;
            if(penultimate_operation = '1') then
                next_state <= square_direct_7;
            end if;
        when square_direct_7 => 
            next_state <= square_direct_7;
            if(penultimate_operation = '1') then
                if(operands_size = "10") then
                    next_state <= square_direct_8;
                else
                    next_state <= square_direct_12;
                end if;
            end if;
        when square_direct_8 => 
            next_state <= square_direct_8;
            if(penultimate_operation = '1') then
                next_state <= square_direct_9;
            end if;
        when square_direct_9 => 
            next_state <= square_direct_9;
            if(penultimate_operation = '1') then
                next_state <= square_direct_10;
            end if;
        when square_direct_10 => 
            next_state <= square_direct_10;
            if(penultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when square_direct_12 => 
            next_state <= square_direct_12;
            if(penultimate_operation = '1') then
                next_state <= square_direct_13;
            end if;
        when square_direct_13 => 
            next_state <= square_direct_13;
            if(penultimate_operation = '1') then
                next_state <= square_direct_14;
            end if;
        when square_direct_14 => 
            next_state <= square_direct_14;
            if(penultimate_operation = '1') then
                next_state <= square_direct_15;
            end if;
        when square_direct_15 => 
            next_state <= square_direct_15;
            if(penultimate_operation = '1') then
                next_state <= square_direct_16;
            end if;
        when square_direct_16 => 
            next_state <= square_direct_16;
            if(penultimate_operation = '1') then
                next_state <= square_direct_17;
            end if;
        when square_direct_17 => 
            next_state <= square_direct_17;
            if(penultimate_operation = '1') then
                next_state <= square_direct_18;
            end if;
        when square_direct_18 => 
            next_state <= square_direct_18;
            if(penultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when multiplication_with_reduction_0 => 
            next_state <= multiplication_with_reduction_0;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_1;
            end if;
        when multiplication_with_reduction_1 => 
            next_state <= multiplication_with_reduction_1;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_2;
            end if;
        when multiplication_with_reduction_2 => 
            next_state <= multiplication_with_reduction_2;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_3;
            end if;
        when multiplication_with_reduction_3 => 
            next_state <= multiplication_with_reduction_3;
            if(penultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when multiplication_with_reduction_5 => 
            next_state <= multiplication_with_reduction_5;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_6;
            end if;
        when multiplication_with_reduction_6 => 
            next_state <= multiplication_with_reduction_6;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_7;
            end if;
        when multiplication_with_reduction_7 => 
            next_state <= multiplication_with_reduction_7;
            if(penultimate_operation = '1') then
                if(operands_size = "01") then
                    next_state <= multiplication_with_reduction_8;
                else
                    next_state <= multiplication_with_reduction_16;
                end if;
            end if;
        when multiplication_with_reduction_8 => 
            next_state <= multiplication_with_reduction_8;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_9;
            end if;
        when multiplication_with_reduction_9 => 
            next_state <= multiplication_with_reduction_9;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_10;
            end if;
        when multiplication_with_reduction_10 => 
            next_state <= multiplication_with_reduction_10;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_11;
            end if;
        when multiplication_with_reduction_11 => 
            next_state <= multiplication_with_reduction_11;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_12;
            end if;
        when multiplication_with_reduction_12 => 
            next_state <= multiplication_with_reduction_12;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_13;
            end if;
        when multiplication_with_reduction_13 => 
            next_state <= multiplication_with_reduction_13;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_14;
            end if;
        when multiplication_with_reduction_14 => 
            next_state <= multiplication_with_reduction_14;
            if(penultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when multiplication_with_reduction_16 => 
            next_state <= multiplication_with_reduction_16;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_17;
            end if;
        when multiplication_with_reduction_17 => 
            next_state <= multiplication_with_reduction_17;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_18;
            end if;
        when multiplication_with_reduction_18 => 
            next_state <= multiplication_with_reduction_18;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_19;
            end if;
        when multiplication_with_reduction_19 => 
            next_state <= multiplication_with_reduction_19;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_20;
            end if;
        when multiplication_with_reduction_20 => 
            next_state <= multiplication_with_reduction_20;
            if(penultimate_operation = '1') then
                if(operands_size = "10") then
                    next_state <= multiplication_with_reduction_21;
                else
                    next_state <= multiplication_with_reduction_35;
                end if;
            end if;
        when multiplication_with_reduction_21 => 
            next_state <= multiplication_with_reduction_21;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_22;
            end if;
        when multiplication_with_reduction_22 => 
            next_state <= multiplication_with_reduction_22;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_23;
            end if;
        when multiplication_with_reduction_23 => 
            next_state <= multiplication_with_reduction_23;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_24;
            end if;
        when multiplication_with_reduction_24 => 
            next_state <= multiplication_with_reduction_24;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_25;
            end if;
        when multiplication_with_reduction_25 => 
            next_state <= multiplication_with_reduction_25;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_26;
            end if;
        when multiplication_with_reduction_26 => 
            next_state <= multiplication_with_reduction_26;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_27;
            end if;
        when multiplication_with_reduction_27 => 
            next_state <= multiplication_with_reduction_27;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_28;
            end if;
        when multiplication_with_reduction_28 => 
            next_state <= multiplication_with_reduction_28;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_29;
            end if;
        when multiplication_with_reduction_29 => 
            next_state <= multiplication_with_reduction_29;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_30;
            end if;
        when multiplication_with_reduction_30 => 
            next_state <= multiplication_with_reduction_30;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_31;
            end if;
        when multiplication_with_reduction_31 => 
            next_state <= multiplication_with_reduction_31;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_32;
            end if;
        when multiplication_with_reduction_32 => 
            next_state <= multiplication_with_reduction_32;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_33;
            end if;
        when multiplication_with_reduction_33 => 
            next_state <= multiplication_with_reduction_33;
            if(penultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
       when multiplication_with_reduction_35 => 
            next_state <= multiplication_with_reduction_35;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_36;
            end if;
        when multiplication_with_reduction_36 => 
            next_state <= multiplication_with_reduction_36;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_37;
            end if;
        when multiplication_with_reduction_37 => 
            next_state <= multiplication_with_reduction_37;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_38;
            end if;
        when multiplication_with_reduction_38 => 
            next_state <= multiplication_with_reduction_38;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_39;
            end if;
        when multiplication_with_reduction_39 => 
            next_state <= multiplication_with_reduction_39;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_40;
            end if;
        when multiplication_with_reduction_40 => 
            next_state <= multiplication_with_reduction_40;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_41;
            end if;
        when multiplication_with_reduction_41 => 
            next_state <= multiplication_with_reduction_41;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_42;
            end if;
        when multiplication_with_reduction_42 => 
            next_state <= multiplication_with_reduction_42;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_43;
            end if;
        when multiplication_with_reduction_43 => 
            next_state <= multiplication_with_reduction_43;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_44;
            end if;
        when multiplication_with_reduction_44 => 
            next_state <= multiplication_with_reduction_44;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_45;
            end if;
        when multiplication_with_reduction_45 => 
            next_state <= multiplication_with_reduction_45;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_46;
            end if;
        when multiplication_with_reduction_46 => 
            next_state <= multiplication_with_reduction_46;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_47;
            end if;
        when multiplication_with_reduction_47 => 
            next_state <= multiplication_with_reduction_47;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_48;
            end if;
        when multiplication_with_reduction_48 => 
            next_state <= multiplication_with_reduction_48;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_49;
            end if;
        when multiplication_with_reduction_49 => 
            next_state <= multiplication_with_reduction_49;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_50;
            end if;
        when multiplication_with_reduction_50 => 
            next_state <= multiplication_with_reduction_50;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_51;
            end if;
        when multiplication_with_reduction_51 => 
            next_state <= multiplication_with_reduction_51;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_52;
            end if;
        when multiplication_with_reduction_52 => 
            next_state <= multiplication_with_reduction_52;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_53;
            end if;
        when multiplication_with_reduction_53 => 
            next_state <= multiplication_with_reduction_53;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_54;
            end if;
        when multiplication_with_reduction_54 => 
            next_state <= multiplication_with_reduction_54;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_55;
            end if;
        when multiplication_with_reduction_55 => 
            next_state <= multiplication_with_reduction_55;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_56;
            end if;
        when multiplication_with_reduction_56 => 
            next_state <= multiplication_with_reduction_56;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_57;
            end if;
        when multiplication_with_reduction_57 => 
            next_state <= multiplication_with_reduction_57;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_58;
            end if;
        when multiplication_with_reduction_58 => 
            next_state <= multiplication_with_reduction_58;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_59;
            end if;
        when multiplication_with_reduction_59 => 
            next_state <= multiplication_with_reduction_59;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_60;
            end if;
        when multiplication_with_reduction_60 => 
            next_state <= multiplication_with_reduction_60;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_61;
            end if;
        when multiplication_with_reduction_61 => 
            next_state <= multiplication_with_reduction_61;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_62;
            end if;
        when multiplication_with_reduction_62 => 
            next_state <= multiplication_with_reduction_62;
            if(penultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when multiplication_with_reduction_special_prime_0 => 
            next_state <= multiplication_with_reduction_special_prime_0;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_1;
            end if;
        when multiplication_with_reduction_special_prime_1 => 
            next_state <= multiplication_with_reduction_special_prime_1;
            if(penultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when multiplication_with_reduction_special_prime_3 => 
            next_state <= multiplication_with_reduction_special_prime_3;
            if(penultimate_operation = '1') then
                if(operands_size = "01") then
                    next_state <= multiplication_with_reduction_special_prime_4;
                else
                    next_state <= multiplication_with_reduction_special_prime_10;
                end if;
            end if;
        when multiplication_with_reduction_special_prime_4 => 
            next_state <= multiplication_with_reduction_special_prime_4;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_5;
            end if;
        when multiplication_with_reduction_special_prime_5 => 
            next_state <= multiplication_with_reduction_special_prime_5;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_6;
            end if;
        when multiplication_with_reduction_special_prime_6 => 
            next_state <= multiplication_with_reduction_special_prime_6;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_7;
            end if;
        when multiplication_with_reduction_special_prime_7 => 
            next_state <= multiplication_with_reduction_special_prime_7;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_8;
            end if;
        when multiplication_with_reduction_special_prime_8 => 
            next_state <= multiplication_with_reduction_special_prime_8;
            if(penultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when multiplication_with_reduction_special_prime_10 => 
            next_state <= multiplication_with_reduction_special_prime_10;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_11;
            end if;
        when multiplication_with_reduction_special_prime_11 => 
            next_state <= multiplication_with_reduction_special_prime_11;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_12;
            end if;
        when multiplication_with_reduction_special_prime_12 => 
            next_state <= multiplication_with_reduction_special_prime_12;
            if(penultimate_operation = '1') then
                if(operands_size = "10") then
                    next_state <= multiplication_with_reduction_special_prime_13;
                else
                    next_state <= multiplication_with_reduction_special_prime_25;
                end if;
            end if;
        when multiplication_with_reduction_special_prime_13 => 
            next_state <= multiplication_with_reduction_special_prime_13;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_14;
            end if;
        when multiplication_with_reduction_special_prime_14 => 
            next_state <= multiplication_with_reduction_special_prime_14;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_15;
            end if;
        when multiplication_with_reduction_special_prime_15 => 
            next_state <= multiplication_with_reduction_special_prime_15;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_16;
            end if;
        when multiplication_with_reduction_special_prime_16 => 
            next_state <= multiplication_with_reduction_special_prime_16;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_17;
            end if;
        when multiplication_with_reduction_special_prime_17 => 
            next_state <= multiplication_with_reduction_special_prime_17;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_18;
            end if;
        when multiplication_with_reduction_special_prime_18 => 
            next_state <= multiplication_with_reduction_special_prime_18;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_19;
            end if;
        when multiplication_with_reduction_special_prime_19 => 
            next_state <= multiplication_with_reduction_special_prime_19;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_20;
            end if;
        when multiplication_with_reduction_special_prime_20 => 
            next_state <= multiplication_with_reduction_special_prime_20;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_21;
            end if;
        when multiplication_with_reduction_special_prime_21 => 
            next_state <= multiplication_with_reduction_special_prime_21;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_22;
            end if;
        when multiplication_with_reduction_special_prime_22 => 
            next_state <= multiplication_with_reduction_special_prime_22;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_23;
            end if;
        when multiplication_with_reduction_special_prime_23 => 
            next_state <= multiplication_with_reduction_special_prime_23;
            if(penultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when multiplication_with_reduction_special_prime_25 => 
            next_state <= multiplication_with_reduction_special_prime_25;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_26;
            end if;
        when multiplication_with_reduction_special_prime_26 => 
            next_state <= multiplication_with_reduction_special_prime_26;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_27;
            end if;
        when multiplication_with_reduction_special_prime_27 => 
            next_state <= multiplication_with_reduction_special_prime_27;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_28;
            end if;
        when multiplication_with_reduction_special_prime_28 => 
            next_state <= multiplication_with_reduction_special_prime_28;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_29;
            end if;
        when multiplication_with_reduction_special_prime_29 => 
            next_state <= multiplication_with_reduction_special_prime_29;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_30;
            end if;
        when multiplication_with_reduction_special_prime_30 => 
            next_state <= multiplication_with_reduction_special_prime_30;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_31;
            end if;
        when multiplication_with_reduction_special_prime_31 => 
            next_state <= multiplication_with_reduction_special_prime_31;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_32;
            end if;
        when multiplication_with_reduction_special_prime_32 => 
            next_state <= multiplication_with_reduction_special_prime_32;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_33;
            end if;
        when multiplication_with_reduction_special_prime_33 => 
            next_state <= multiplication_with_reduction_special_prime_33;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_34;
            end if;
        when multiplication_with_reduction_special_prime_34 => 
            next_state <= multiplication_with_reduction_special_prime_34;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_35;
            end if;
        when multiplication_with_reduction_special_prime_35 => 
            next_state <= multiplication_with_reduction_special_prime_35;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_36;
            end if;
        when multiplication_with_reduction_special_prime_36 => 
            next_state <= multiplication_with_reduction_special_prime_36;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_37;
            end if;
        when multiplication_with_reduction_special_prime_37 => 
            next_state <= multiplication_with_reduction_special_prime_37;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_38;
            end if;
        when multiplication_with_reduction_special_prime_38 => 
            next_state <= multiplication_with_reduction_special_prime_38;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_39;
            end if;
        when multiplication_with_reduction_special_prime_39 => 
            next_state <= multiplication_with_reduction_special_prime_39;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_40;
            end if;
        when multiplication_with_reduction_special_prime_40 => 
            next_state <= multiplication_with_reduction_special_prime_40;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_41;
            end if;
        when multiplication_with_reduction_special_prime_41 => 
            next_state <= multiplication_with_reduction_special_prime_41;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_42;
            end if;
        when multiplication_with_reduction_special_prime_42 => 
            next_state <= multiplication_with_reduction_special_prime_42;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_43;
            end if;
        when multiplication_with_reduction_special_prime_43 => 
            next_state <= multiplication_with_reduction_special_prime_43;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_44;
            end if;
        when multiplication_with_reduction_special_prime_44 => 
            next_state <= multiplication_with_reduction_special_prime_44;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_45;
            end if;
        when multiplication_with_reduction_special_prime_45 => 
            next_state <= multiplication_with_reduction_special_prime_45;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_46;
            end if;
        when multiplication_with_reduction_special_prime_46 => 
            next_state <= multiplication_with_reduction_special_prime_46;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_47;
            end if;
        when multiplication_with_reduction_special_prime_47 => 
            next_state <= multiplication_with_reduction_special_prime_47;
            if(penultimate_operation = '1') then
                next_state <= multiplication_with_reduction_special_prime_48;
            end if;
        when multiplication_with_reduction_special_prime_48 => 
            next_state <= multiplication_with_reduction_special_prime_48;
            if(penultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when square_with_reduction_0 => 
            next_state <= square_with_reduction_0;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_1;
            end if;
        when square_with_reduction_1 => 
            next_state <= square_with_reduction_1;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_2;
            end if;
        when square_with_reduction_2 => 
            next_state <= square_with_reduction_2;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_3;
            end if;
        when square_with_reduction_3 => 
            next_state <= square_with_reduction_3;
            if(penultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when square_with_reduction_5 => 
            next_state <= square_with_reduction_5;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_6;
            end if;
        when square_with_reduction_6 => 
            next_state <= square_with_reduction_6;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_7;
            end if;
        when square_with_reduction_7 => 
            next_state <= square_with_reduction_7;
            if(penultimate_operation = '1') then
                if(operands_size = "01") then
                    next_state <= square_with_reduction_8;
                else
                    next_state <= square_with_reduction_15;
                end if;
            end if;
        when square_with_reduction_8 => 
            next_state <= square_with_reduction_8;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_9;
            end if;
        when square_with_reduction_9 => 
            next_state <= square_with_reduction_9;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_10;
            end if;
        when square_with_reduction_10 => 
            next_state <= square_with_reduction_10;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_11;
            end if;
        when square_with_reduction_11 => 
            next_state <= square_with_reduction_11;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_12;
            end if;
        when square_with_reduction_12 => 
            next_state <= square_with_reduction_12;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_13;
            end if;
        when square_with_reduction_13 => 
            next_state <= square_with_reduction_13;
            if(penultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when square_with_reduction_15 => 
            next_state <= square_with_reduction_15;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_16;
            end if;
        when square_with_reduction_16 => 
            next_state <= square_with_reduction_16;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_17;
            end if;
        when square_with_reduction_17 => 
            next_state <= square_with_reduction_17;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_18;
            end if;
        when square_with_reduction_18 => 
            next_state <= square_with_reduction_18;
            if(penultimate_operation = '1') then
                if(operands_size = "10") then
                    next_state <= square_with_reduction_19;
                else
                    next_state <= square_with_reduction_31;
                end if;
            end if;
        when square_with_reduction_19 => 
            next_state <= square_with_reduction_19;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_20;
            end if;
        when square_with_reduction_20 => 
            next_state <= square_with_reduction_20;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_21;
            end if;
        when square_with_reduction_21 => 
            next_state <= square_with_reduction_21;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_22;
            end if;
        when square_with_reduction_22 => 
            next_state <= square_with_reduction_22;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_23;
            end if;
        when square_with_reduction_23 => 
            next_state <= square_with_reduction_23;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_24;
            end if;
        when square_with_reduction_24 => 
            next_state <= square_with_reduction_24;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_25;
            end if;
        when square_with_reduction_25 => 
            next_state <= square_with_reduction_25;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_26;
            end if;
        when square_with_reduction_26 => 
            next_state <= square_with_reduction_26;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_27;
            end if;
        when square_with_reduction_27 => 
            next_state <= square_with_reduction_27;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_28;
            end if;
        when square_with_reduction_28 => 
            next_state <= square_with_reduction_28;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_29;
            end if;
        when square_with_reduction_29 => 
            next_state <= square_with_reduction_29;
            if(penultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when square_with_reduction_31 => 
            next_state <= square_with_reduction_31;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_32;
            end if;
        when square_with_reduction_32 => 
            next_state <= square_with_reduction_32;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_33;
            end if;
        when square_with_reduction_33 => 
            next_state <= square_with_reduction_33;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_34;
            end if;
        when square_with_reduction_34 => 
            next_state <= square_with_reduction_34;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_35;
            end if;
        when square_with_reduction_35 => 
            next_state <= square_with_reduction_35;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_36;
            end if;
        when square_with_reduction_36 => 
            next_state <= square_with_reduction_36;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_37;
            end if;
        when square_with_reduction_37 => 
            next_state <= square_with_reduction_37;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_38;
            end if;
        when square_with_reduction_38 => 
            next_state <= square_with_reduction_38;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_39;
            end if;
        when square_with_reduction_39 => 
            next_state <= square_with_reduction_39;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_40;
            end if;
        when square_with_reduction_40 => 
            next_state <= square_with_reduction_40;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_41;
            end if;
        when square_with_reduction_41 => 
            next_state <= square_with_reduction_41;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_42;
            end if;
        when square_with_reduction_42 => 
            next_state <= square_with_reduction_42;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_43;
            end if;
        when square_with_reduction_43 => 
            next_state <= square_with_reduction_43;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_44;
            end if;
        when square_with_reduction_44 => 
            next_state <= square_with_reduction_44;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_45;
            end if;
        when square_with_reduction_45 => 
            next_state <= square_with_reduction_45;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_46;
            end if;
        when square_with_reduction_46 => 
            next_state <= square_with_reduction_46;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_47;
            end if;
        when square_with_reduction_47 => 
            next_state <= square_with_reduction_47;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_48;
            end if;
        when square_with_reduction_48 => 
            next_state <= square_with_reduction_48;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_49;
            end if;
        when square_with_reduction_49 => 
            next_state <= square_with_reduction_49;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_50;
            end if;
        when square_with_reduction_50 => 
            next_state <= square_with_reduction_50;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_51;
            end if;
        when square_with_reduction_51 => 
            next_state <= square_with_reduction_51;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_52;
            end if;
        when square_with_reduction_52 => 
            next_state <= square_with_reduction_52;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_53;
            end if;
        when square_with_reduction_53 => 
            next_state <= square_with_reduction_53;
            if(penultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when square_with_reduction_special_prime_0 => 
            next_state <= square_with_reduction_special_prime_0;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_1;
            end if;
        when square_with_reduction_special_prime_1 => 
            next_state <= square_with_reduction_special_prime_1;
            if(penultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when square_with_reduction_special_prime_3 => 
            next_state <= square_with_reduction_special_prime_3;
            if(penultimate_operation = '1') then
                if(operands_size = "01") then
                    next_state <= square_with_reduction_special_prime_4;
                else
                    next_state <= square_with_reduction_special_prime_9;
                end if;
            end if;
        when square_with_reduction_special_prime_4 =>
            next_state <= square_with_reduction_special_prime_4;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_5;
            end if;
        when square_with_reduction_special_prime_5 => 
            next_state <= square_with_reduction_special_prime_5;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_6;
            end if;
        when square_with_reduction_special_prime_6 => 
            next_state <= square_with_reduction_special_prime_6;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_7;
            end if;
        when square_with_reduction_special_prime_7 => 
            next_state <= square_with_reduction_special_prime_7;
            if(penultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when square_with_reduction_special_prime_9 => 
            next_state <= square_with_reduction_special_prime_9;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_10;
            end if;
        when square_with_reduction_special_prime_10 => 
            next_state <= square_with_reduction_special_prime_10;
            if(penultimate_operation = '1') then
                if(operands_size = "10") then
                    next_state <= square_with_reduction_special_prime_11;
                else
                    next_state <= square_with_reduction_special_prime_21;
                end if;
            end if;
        when square_with_reduction_special_prime_11 => 
            next_state <= square_with_reduction_special_prime_11;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_12;
            end if;
        when square_with_reduction_special_prime_12 => 
            next_state <= square_with_reduction_special_prime_12;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_13;
            end if;
        when square_with_reduction_special_prime_13 => 
            next_state <= square_with_reduction_special_prime_13;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_14;
            end if;
        when square_with_reduction_special_prime_14 => 
            next_state <= square_with_reduction_special_prime_14;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_15;
            end if;
        when square_with_reduction_special_prime_15 => 
            next_state <= square_with_reduction_special_prime_15;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_16;
            end if;
        when square_with_reduction_special_prime_16 => 
            next_state <= square_with_reduction_special_prime_16;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_17;
            end if;
        when square_with_reduction_special_prime_17 => 
            next_state <= square_with_reduction_special_prime_17;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_18;
            end if;
        when square_with_reduction_special_prime_18 => 
            next_state <= square_with_reduction_special_prime_18;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_19;
            end if;
        when square_with_reduction_special_prime_19 => 
            next_state <= square_with_reduction_special_prime_19;
            if(penultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
        when square_with_reduction_special_prime_21 => 
            next_state <= square_with_reduction_special_prime_21;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_22;
            end if;
        when square_with_reduction_special_prime_22 => 
            next_state <= square_with_reduction_special_prime_22;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_23;
            end if;
        when square_with_reduction_special_prime_23 => 
            next_state <= square_with_reduction_special_prime_23;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_24;
            end if;
        when square_with_reduction_special_prime_24 => 
            next_state <= square_with_reduction_special_prime_24;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_25;
            end if;
        when square_with_reduction_special_prime_25 => 
            next_state <= square_with_reduction_special_prime_25;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_26;
            end if;
        when square_with_reduction_special_prime_26 => 
            next_state <= square_with_reduction_special_prime_26;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_27;
            end if;
        when square_with_reduction_special_prime_27 => 
            next_state <= square_with_reduction_special_prime_27;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_28;
            end if;
        when square_with_reduction_special_prime_28 => 
            next_state <= square_with_reduction_special_prime_28;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_29;
            end if;
        when square_with_reduction_special_prime_29 => 
            next_state <= square_with_reduction_special_prime_29;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_30;
            end if;
        when square_with_reduction_special_prime_30 => 
            next_state <= square_with_reduction_special_prime_30;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_31;
            end if;
        when square_with_reduction_special_prime_31 => 
            next_state <= square_with_reduction_special_prime_31;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_32;
            end if;
        when square_with_reduction_special_prime_32 => 
            next_state <= square_with_reduction_special_prime_32;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_33;
            end if;
        when square_with_reduction_special_prime_33 => 
            next_state <= square_with_reduction_special_prime_33;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_34;
            end if;
        when square_with_reduction_special_prime_34 => 
            next_state <= square_with_reduction_special_prime_34;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_35;
            end if;
        when square_with_reduction_special_prime_35 => 
            next_state <= square_with_reduction_special_prime_35;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_36;
            end if;
        when square_with_reduction_special_prime_36 => 
            next_state <= square_with_reduction_special_prime_36;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_37;
            end if;
        when square_with_reduction_special_prime_37 => 
            next_state <= square_with_reduction_special_prime_37;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_38;
            end if;
        when square_with_reduction_special_prime_38 => 
            next_state <= square_with_reduction_special_prime_38;
            if(penultimate_operation = '1') then
                next_state <= square_with_reduction_special_prime_39;
            end if;
        when square_with_reduction_special_prime_39 => 
            next_state <= square_with_reduction_special_prime_39;
            if(penultimate_operation = '1') then
                next_state <= nop_8_stages;
            end if;
            
        when addition_subtraction_direct_0 =>
            next_state <= addition_subtraction_direct_0;
            if(penultimate_operation = '1') then
                next_state <= nop_4_stages;
            end if;
        when addition_subtraction_direct_2 =>
            next_state <= addition_subtraction_direct_2;
            if(penultimate_operation = '1') then
                if(operands_size = "01") then
                    next_state <= addition_subtraction_direct_3;
                else
                    next_state <= addition_subtraction_direct_5;
                end if;
            end if;
        when addition_subtraction_direct_3 =>
            next_state <= addition_subtraction_direct_3;
            if(penultimate_operation = '1') then
                next_state <= nop_4_stages;
            end if;
        when addition_subtraction_direct_5 =>
            next_state <= addition_subtraction_direct_5;
            if(penultimate_operation = '1') then
                if(operands_size = "10") then
                    next_state <= addition_subtraction_direct_6;
                else
                    next_state <= addition_subtraction_direct_8;
                end if;
            end if;
        when addition_subtraction_direct_6 =>
            next_state <= addition_subtraction_direct_6;
            if(penultimate_operation = '1') then
                next_state <= nop_4_stages;
            end if;
        when addition_subtraction_direct_8 =>
            next_state <= addition_subtraction_direct_8;
            if(penultimate_operation = '1') then
                next_state <= addition_subtraction_direct_9;
            end if;
        when addition_subtraction_direct_9 =>
            next_state <= addition_subtraction_direct_9;
            if(penultimate_operation = '1') then
                next_state <= nop_4_stages;
            end if;
        when iterative_modular_reduction_0 =>
            next_state <= iterative_modular_reduction_0;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_1;
            end if;    
        when iterative_modular_reduction_1 =>
            next_state <= iterative_modular_reduction_1;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_2;
            end if;
        when iterative_modular_reduction_2 =>
            next_state <= iterative_modular_reduction_2;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_3;
            end if;
        when iterative_modular_reduction_3 =>
            next_state <= iterative_modular_reduction_3;
            if(penultimate_operation = '1') then
                next_state <= nop_4_stages;
            end if;
        when iterative_modular_reduction_5 =>
            next_state <= iterative_modular_reduction_5;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_6;
            end if;
        when iterative_modular_reduction_6 =>
            next_state <= iterative_modular_reduction_6;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_7;
            end if;
        when iterative_modular_reduction_7 =>
            next_state <= iterative_modular_reduction_7;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_8;
            end if;
        when iterative_modular_reduction_8 =>
            next_state <= iterative_modular_reduction_8;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_9;
            end if;
        when iterative_modular_reduction_9 =>
            next_state <= iterative_modular_reduction_9;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_10;
            end if;
        when iterative_modular_reduction_10 =>
            next_state <= iterative_modular_reduction_10;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_11;
            end if;
        when iterative_modular_reduction_11 =>
            next_state <= iterative_modular_reduction_11;
            if(penultimate_operation = '1') then
                next_state <= nop_4_stages;
            end if;
        when iterative_modular_reduction_13 =>
            next_state <= iterative_modular_reduction_13;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_14;
            end if;
        when iterative_modular_reduction_14 =>
            next_state <= iterative_modular_reduction_14;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_15;
            end if;
        when iterative_modular_reduction_15 =>
            next_state <= iterative_modular_reduction_15;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_16;
            end if;
        when iterative_modular_reduction_16 =>
            next_state <= iterative_modular_reduction_16;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_17;
            end if;
        when iterative_modular_reduction_17 =>
            next_state <= iterative_modular_reduction_17;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_18;
            end if;
        when iterative_modular_reduction_18 =>
            next_state <= iterative_modular_reduction_18;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_19;
            end if;
        when iterative_modular_reduction_19 =>
            next_state <= iterative_modular_reduction_19;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_20;
            end if;
        when iterative_modular_reduction_20 =>
            next_state <= iterative_modular_reduction_20;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_21;
            end if;
        when iterative_modular_reduction_21 =>
            next_state <= iterative_modular_reduction_21;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_22;
            end if;
        when iterative_modular_reduction_22 =>
            next_state <= iterative_modular_reduction_22;
            if(penultimate_operation = '1') then
                next_state <= nop_4_stages;
            end if;
        when iterative_modular_reduction_24 =>
            next_state <= iterative_modular_reduction_24;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_25;
            end if;
        when iterative_modular_reduction_25 =>
            next_state <= iterative_modular_reduction_25;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_26;
            end if;
        when iterative_modular_reduction_26 =>
            next_state <= iterative_modular_reduction_26;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_27;
            end if;
        when iterative_modular_reduction_27 =>
            next_state <= iterative_modular_reduction_27;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_28;
            end if;
        when iterative_modular_reduction_28 =>
            next_state <= iterative_modular_reduction_28;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_29;
            end if;
        when iterative_modular_reduction_29 =>
            next_state <= iterative_modular_reduction_29;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_30;
            end if;
        when iterative_modular_reduction_30 =>
            next_state <= iterative_modular_reduction_30;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_31;
            end if;
        when iterative_modular_reduction_31 =>
            next_state <= iterative_modular_reduction_31;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_32;
            end if;
        when iterative_modular_reduction_32 =>
            next_state <= iterative_modular_reduction_32;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_33;
            end if;
        when iterative_modular_reduction_33 =>
            next_state <= iterative_modular_reduction_33;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_34;
            end if;
        when iterative_modular_reduction_34 =>
            next_state <= iterative_modular_reduction_34;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_35;
            end if;
        when iterative_modular_reduction_35 =>
            next_state <= iterative_modular_reduction_35;
            if(penultimate_operation = '1') then
                next_state <= iterative_modular_reduction_36;
            end if;
        when iterative_modular_reduction_36 =>
            next_state <= iterative_modular_reduction_36;
            if(penultimate_operation = '1') then
                next_state <= nop_4_stages;
            end if;
        when nop_4_stages =>
            next_state <= nop_4_stages;
            if(penultimate_operation = '1') then
                next_state <= decode_instruction;
            end if;
        when nop_8_stages =>
            next_state <= nop_8_stages;
            if(penultimate_operation = '1') then
                next_state <= decode_instruction;
            end if;
    end case;
end process;

end behavioral;