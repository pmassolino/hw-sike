----------------------------------------------------------------------------------
-- Implementation by Pedro Maat C. Massolino,
-- hereby denoted as "the implementer".
--
-- To the extent possible under law, the implementer has waived all copyright
-- and related or neighboring rights to the source code in this file.
-- http://creativecommons.org/publicdomain/zero/1.0/
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

architecture tiled_behavioral_v1 of pipeline_signed_base_multiplier_257 is

signal temp_mult_0 : std_logic_vector(40 downto 0);
signal temp_mult_1 : std_logic_vector(64 downto 24);
signal temp_mult_2 : std_logic_vector(88 downto 48);
signal temp_mult_3 : std_logic_vector(112 downto 72);
signal temp_mult_4 : std_logic_vector(136 downto 96);
signal temp_mult_5 : std_logic_vector(57 downto 17);
signal temp_mult_6 : std_logic_vector(81 downto 41);
signal temp_mult_7 : std_logic_vector(105 downto 65);
signal temp_mult_8 : std_logic_vector(129 downto 89);
signal temp_mult_9 : std_logic_vector(153 downto 113);
signal temp_mult_10 : std_logic_vector(74 downto 34);
signal temp_mult_11 : std_logic_vector(98 downto 58);
signal temp_mult_12 : std_logic_vector(122 downto 82);
signal temp_mult_13 : std_logic_vector(146 downto 106);
signal temp_mult_14 : std_logic_vector(170 downto 130);
signal temp_mult_15 : std_logic_vector(91 downto 51);
signal temp_mult_16 : std_logic_vector(115 downto 75);
signal temp_mult_17 : std_logic_vector(139 downto 99);
signal temp_mult_18 : std_logic_vector(163 downto 123);
signal temp_mult_19 : std_logic_vector(187 downto 147);
signal temp_mult_20 : std_logic_vector(108 downto 68);
signal temp_mult_21 : std_logic_vector(132 downto 92);
signal temp_mult_22 : std_logic_vector(156 downto 116);
signal temp_mult_23 : std_logic_vector(180 downto 140);
signal temp_mult_24 : std_logic_vector(204 downto 164);
signal temp_mult_25 : std_logic_vector(125 downto 85);
signal temp_mult_26 : std_logic_vector(149 downto 109);
signal temp_mult_27 : std_logic_vector(173 downto 133);
signal temp_mult_28 : std_logic_vector(197 downto 157);
signal temp_mult_29 : std_logic_vector(221 downto 181);
signal temp_mult_30 : std_logic_vector(142 downto 102);
signal temp_mult_31 : std_logic_vector(166 downto 126);
signal temp_mult_32 : std_logic_vector(190 downto 150);
signal temp_mult_33 : std_logic_vector(214 downto 174);
signal temp_mult_34 : std_logic_vector(238 downto 198);
signal temp_mult_35 : std_logic_vector(159 downto 119);
signal temp_mult_36 : std_logic_vector(183 downto 143);
signal temp_mult_37 : std_logic_vector(207 downto 167);
signal temp_mult_38 : std_logic_vector(231 downto 191);
signal temp_mult_39 : std_logic_vector(255 downto 215);
signal temp_mult_40 : std_logic_vector(160 downto 120);
signal temp_mult_41 : std_logic_vector(177 downto 137);
signal temp_mult_42 : std_logic_vector(194 downto 154);
signal temp_mult_43 : std_logic_vector(211 downto 171);
signal temp_mult_44 : std_logic_vector(228 downto 188);
signal temp_mult_45 : std_logic_vector(245 downto 205);
signal temp_mult_46 : std_logic_vector(262 downto 222);
signal temp_mult_47 : std_logic_vector(279 downto 239);
signal temp_mult_48 : std_logic_vector(184 downto 144);
signal temp_mult_49 : std_logic_vector(201 downto 161);
signal temp_mult_50 : std_logic_vector(218 downto 178);
signal temp_mult_51 : std_logic_vector(235 downto 195);
signal temp_mult_52 : std_logic_vector(252 downto 212);
signal temp_mult_53 : std_logic_vector(269 downto 229);
signal temp_mult_54 : std_logic_vector(286 downto 246);
signal temp_mult_55 : std_logic_vector(303 downto 263);
signal temp_mult_56 : std_logic_vector(208 downto 168);
signal temp_mult_57 : std_logic_vector(225 downto 185);
signal temp_mult_58 : std_logic_vector(242 downto 202);
signal temp_mult_59 : std_logic_vector(259 downto 219);
signal temp_mult_60 : std_logic_vector(276 downto 236);
signal temp_mult_61 : std_logic_vector(293 downto 253);
signal temp_mult_62 : std_logic_vector(310 downto 270);
signal temp_mult_63 : std_logic_vector(327 downto 287);
signal temp_mult_64 : std_logic_vector(232 downto 192);
signal temp_mult_65 : std_logic_vector(249 downto 209);
signal temp_mult_66 : std_logic_vector(266 downto 226);
signal temp_mult_67 : std_logic_vector(283 downto 243);
signal temp_mult_68 : std_logic_vector(300 downto 260);
signal temp_mult_69 : std_logic_vector(317 downto 277);
signal temp_mult_70 : std_logic_vector(334 downto 294);
signal temp_mult_71 : std_logic_vector(351 downto 311);
signal temp_mult_72 : std_logic_vector(256 downto 216);
signal temp_mult_73 : std_logic_vector(273 downto 233);
signal temp_mult_74 : std_logic_vector(290 downto 250);
signal temp_mult_75 : std_logic_vector(307 downto 267);
signal temp_mult_76 : std_logic_vector(324 downto 284);
signal temp_mult_77 : std_logic_vector(341 downto 301);
signal temp_mult_78 : std_logic_vector(358 downto 318);
signal temp_mult_79 : std_logic_vector(375 downto 335);
signal temp_mult_80 : std_logic_vector(176 downto 136);
signal temp_mult_81 : std_logic_vector(193 downto 153);
signal temp_mult_82 : std_logic_vector(210 downto 170);
signal temp_mult_83 : std_logic_vector(227 downto 187);
signal temp_mult_84 : std_logic_vector(244 downto 204);
signal temp_mult_85 : std_logic_vector(261 downto 221);
signal temp_mult_86 : std_logic_vector(278 downto 238);
signal temp_mult_87 : std_logic_vector(295 downto 255);
signal temp_mult_88 : std_logic_vector(200 downto 160);
signal temp_mult_89 : std_logic_vector(217 downto 177);
signal temp_mult_90 : std_logic_vector(234 downto 194);
signal temp_mult_91 : std_logic_vector(251 downto 211);
signal temp_mult_92 : std_logic_vector(268 downto 228);
signal temp_mult_93 : std_logic_vector(285 downto 245);
signal temp_mult_94 : std_logic_vector(302 downto 262);
signal temp_mult_95 : std_logic_vector(319 downto 279);
signal temp_mult_96 : std_logic_vector(224 downto 184);
signal temp_mult_97 : std_logic_vector(241 downto 201);
signal temp_mult_98 : std_logic_vector(258 downto 218);
signal temp_mult_99 : std_logic_vector(275 downto 235);
signal temp_mult_100 : std_logic_vector(292 downto 252);
signal temp_mult_101 : std_logic_vector(309 downto 269);
signal temp_mult_102 : std_logic_vector(326 downto 286);
signal temp_mult_103 : std_logic_vector(343 downto 303);
signal temp_mult_104 : std_logic_vector(248 downto 208);
signal temp_mult_105 : std_logic_vector(265 downto 225);
signal temp_mult_106 : std_logic_vector(282 downto 242);
signal temp_mult_107 : std_logic_vector(299 downto 259);
signal temp_mult_108 : std_logic_vector(316 downto 276);
signal temp_mult_109 : std_logic_vector(333 downto 293);
signal temp_mult_110 : std_logic_vector(350 downto 310);
signal temp_mult_111 : std_logic_vector(367 downto 327);
signal temp_mult_112 : std_logic_vector(272 downto 232);
signal temp_mult_113 : std_logic_vector(289 downto 249);
signal temp_mult_114 : std_logic_vector(306 downto 266);
signal temp_mult_115 : std_logic_vector(323 downto 283);
signal temp_mult_116 : std_logic_vector(340 downto 300);
signal temp_mult_117 : std_logic_vector(357 downto 317);
signal temp_mult_118 : std_logic_vector(374 downto 334);
signal temp_mult_119 : std_logic_vector(391 downto 351);
signal temp_mult_120 : std_logic_vector(296 downto 256);
signal temp_mult_121 : std_logic_vector(320 downto 280);
signal temp_mult_122 : std_logic_vector(344 downto 304);
signal temp_mult_123 : std_logic_vector(368 downto 328);
signal temp_mult_124 : std_logic_vector(392 downto 352);
signal temp_mult_125 : std_logic_vector(313 downto 273);
signal temp_mult_126 : std_logic_vector(337 downto 297);
signal temp_mult_127 : std_logic_vector(361 downto 321);
signal temp_mult_128 : std_logic_vector(385 downto 345);
signal temp_mult_129 : std_logic_vector(409 downto 369);
signal temp_mult_130 : std_logic_vector(330 downto 290);
signal temp_mult_131 : std_logic_vector(354 downto 314);
signal temp_mult_132 : std_logic_vector(378 downto 338);
signal temp_mult_133 : std_logic_vector(402 downto 362);
signal temp_mult_134 : std_logic_vector(426 downto 386);
signal temp_mult_135 : std_logic_vector(347 downto 307);
signal temp_mult_136 : std_logic_vector(371 downto 331);
signal temp_mult_137 : std_logic_vector(395 downto 355);
signal temp_mult_138 : std_logic_vector(419 downto 379);
signal temp_mult_139 : std_logic_vector(443 downto 403);
signal temp_mult_140 : std_logic_vector(364 downto 324);
signal temp_mult_141 : std_logic_vector(388 downto 348);
signal temp_mult_142 : std_logic_vector(412 downto 372);
signal temp_mult_143 : std_logic_vector(436 downto 396);
signal temp_mult_144 : std_logic_vector(460 downto 420);
signal temp_mult_145 : std_logic_vector(381 downto 341);
signal temp_mult_146 : std_logic_vector(405 downto 365);
signal temp_mult_147 : std_logic_vector(429 downto 389);
signal temp_mult_148 : std_logic_vector(453 downto 413);
signal temp_mult_149 : std_logic_vector(477 downto 437);
signal temp_mult_150 : std_logic_vector(398 downto 358);
signal temp_mult_151 : std_logic_vector(422 downto 382);
signal temp_mult_152 : std_logic_vector(446 downto 406);
signal temp_mult_153 : std_logic_vector(470 downto 430);
signal temp_mult_154 : std_logic_vector(494 downto 454);
signal temp_mult_155 : std_logic_vector(415 downto 375);
signal temp_mult_156 : std_logic_vector(439 downto 399);
signal temp_mult_157 : std_logic_vector(463 downto 423);
signal temp_mult_158 : std_logic_vector(487 downto 447);
signal temp_mult_159 : std_logic_vector(511 downto 471);
signal temp_mult_160 : std_logic_vector(271 downto 240);
signal temp_part_mult_161 : std_logic_vector(511 downto 256);
signal temp_part_mult_162 : std_logic_vector(512 downto 256);
signal temp_mult_161 : std_logic_vector(513 downto 256);
signal temp_mult_162 : std_logic_vector(513 downto 256);

signal partial_product_0 : std_logic_vector(512 downto 0);
signal partial_product_1 : std_logic_vector(512 downto 0);
signal partial_product_2 : std_logic_vector(512 downto 0);
signal partial_product_3 : std_logic_vector(512 downto 0);
signal partial_product_4 : std_logic_vector(512 downto 0);
signal partial_product_5 : std_logic_vector(512 downto 0);
signal partial_product_6 : std_logic_vector(512 downto 0);
signal partial_product_7 : std_logic_vector(512 downto 0);
signal partial_product_8 : std_logic_vector(512 downto 0);
signal partial_product_9 : std_logic_vector(512 downto 0);
signal partial_product_10 : std_logic_vector(512 downto 0);
signal partial_product_11 : std_logic_vector(512 downto 0);
signal partial_product_12 : std_logic_vector(512 downto 0);
signal partial_product_13 : std_logic_vector(512 downto 0);
signal partial_product_14 : std_logic_vector(512 downto 0);
signal partial_product_15 : std_logic_vector(512 downto 0);
signal partial_product_16 : std_logic_vector(512 downto 0);
signal partial_product_17 : std_logic_vector(512 downto 0);
signal partial_product_18 : std_logic_vector(512 downto 0);
signal partial_product_19 : std_logic_vector(512 downto 0);
signal partial_product_20 : std_logic_vector(512 downto 0);
signal partial_product_21 : std_logic_vector(512 downto 0);
signal partial_product_22 : std_logic_vector(512 downto 0);
signal partial_product_23 : std_logic_vector(512 downto 0);
signal partial_product_24 : std_logic_vector(512 downto 0);
signal partial_product_25 : std_logic_vector(512 downto 0);
signal partial_product_26 : std_logic_vector(513 downto 0);
signal partial_product_27 : std_logic_vector(513 downto 0);

signal temp_o1 : signed(513 downto 0);
signal temp_o2 : signed(513 downto 0);
signal temp_o3 : signed(513 downto 0);
signal temp_o4 : signed(513 downto 0);
signal temp_o5 : signed(513 downto 0);

begin

temp_mult_0 <= std_logic_vector(unsigned(a(16 downto 0)) * unsigned(b(23 downto 0))); 
temp_mult_1 <= std_logic_vector(unsigned(a(16 downto 0)) * unsigned(b(47 downto 24))); 
temp_mult_2 <= std_logic_vector(unsigned(a(16 downto 0)) * unsigned(b(71 downto 48))); 
temp_mult_3 <= std_logic_vector(unsigned(a(16 downto 0)) * unsigned(b(95 downto 72))); 
temp_mult_4 <= std_logic_vector(unsigned(a(16 downto 0)) * unsigned(b(119 downto 96))); 
temp_mult_5 <= std_logic_vector(unsigned(a(33 downto 17)) * unsigned(b(23 downto 0))); 
temp_mult_6 <= std_logic_vector(unsigned(a(33 downto 17)) * unsigned(b(47 downto 24))); 
temp_mult_7 <= std_logic_vector(unsigned(a(33 downto 17)) * unsigned(b(71 downto 48))); 
temp_mult_8 <= std_logic_vector(unsigned(a(33 downto 17)) * unsigned(b(95 downto 72))); 
temp_mult_9 <= std_logic_vector(unsigned(a(33 downto 17)) * unsigned(b(119 downto 96))); 
temp_mult_10 <= std_logic_vector(unsigned(a(50 downto 34)) * unsigned(b(23 downto 0))); 
temp_mult_11 <= std_logic_vector(unsigned(a(50 downto 34)) * unsigned(b(47 downto 24))); 
temp_mult_12 <= std_logic_vector(unsigned(a(50 downto 34)) * unsigned(b(71 downto 48))); 
temp_mult_13 <= std_logic_vector(unsigned(a(50 downto 34)) * unsigned(b(95 downto 72))); 
temp_mult_14 <= std_logic_vector(unsigned(a(50 downto 34)) * unsigned(b(119 downto 96))); 
temp_mult_15 <= std_logic_vector(unsigned(a(67 downto 51)) * unsigned(b(23 downto 0))); 
temp_mult_16 <= std_logic_vector(unsigned(a(67 downto 51)) * unsigned(b(47 downto 24))); 
temp_mult_17 <= std_logic_vector(unsigned(a(67 downto 51)) * unsigned(b(71 downto 48))); 
temp_mult_18 <= std_logic_vector(unsigned(a(67 downto 51)) * unsigned(b(95 downto 72))); 
temp_mult_19 <= std_logic_vector(unsigned(a(67 downto 51)) * unsigned(b(119 downto 96))); 
temp_mult_20 <= std_logic_vector(unsigned(a(84 downto 68)) * unsigned(b(23 downto 0))); 
temp_mult_21 <= std_logic_vector(unsigned(a(84 downto 68)) * unsigned(b(47 downto 24))); 
temp_mult_22 <= std_logic_vector(unsigned(a(84 downto 68)) * unsigned(b(71 downto 48))); 
temp_mult_23 <= std_logic_vector(unsigned(a(84 downto 68)) * unsigned(b(95 downto 72))); 
temp_mult_24 <= std_logic_vector(unsigned(a(84 downto 68)) * unsigned(b(119 downto 96))); 
temp_mult_25 <= std_logic_vector(unsigned(a(101 downto 85)) * unsigned(b(23 downto 0))); 
temp_mult_26 <= std_logic_vector(unsigned(a(101 downto 85)) * unsigned(b(47 downto 24))); 
temp_mult_27 <= std_logic_vector(unsigned(a(101 downto 85)) * unsigned(b(71 downto 48))); 
temp_mult_28 <= std_logic_vector(unsigned(a(101 downto 85)) * unsigned(b(95 downto 72))); 
temp_mult_29 <= std_logic_vector(unsigned(a(101 downto 85)) * unsigned(b(119 downto 96))); 
temp_mult_30 <= std_logic_vector(unsigned(a(118 downto 102)) * unsigned(b(23 downto 0))); 
temp_mult_31 <= std_logic_vector(unsigned(a(118 downto 102)) * unsigned(b(47 downto 24))); 
temp_mult_32 <= std_logic_vector(unsigned(a(118 downto 102)) * unsigned(b(71 downto 48))); 
temp_mult_33 <= std_logic_vector(unsigned(a(118 downto 102)) * unsigned(b(95 downto 72))); 
temp_mult_34 <= std_logic_vector(unsigned(a(118 downto 102)) * unsigned(b(119 downto 96))); 
temp_mult_35 <= std_logic_vector(unsigned(a(135 downto 119)) * unsigned(b(23 downto 0))); 
temp_mult_36 <= std_logic_vector(unsigned(a(135 downto 119)) * unsigned(b(47 downto 24))); 
temp_mult_37 <= std_logic_vector(unsigned(a(135 downto 119)) * unsigned(b(71 downto 48))); 
temp_mult_38 <= std_logic_vector(unsigned(a(135 downto 119)) * unsigned(b(95 downto 72))); 
temp_mult_39 <= std_logic_vector(unsigned(a(135 downto 119)) * unsigned(b(119 downto 96))); 
temp_mult_40 <= std_logic_vector(unsigned(a(23 downto 0)) * unsigned(b(136 downto 120))); 
temp_mult_41 <= std_logic_vector(unsigned(a(23 downto 0)) * unsigned(b(153 downto 137))); 
temp_mult_42 <= std_logic_vector(unsigned(a(23 downto 0)) * unsigned(b(170 downto 154))); 
temp_mult_43 <= std_logic_vector(unsigned(a(23 downto 0)) * unsigned(b(187 downto 171))); 
temp_mult_44 <= std_logic_vector(unsigned(a(23 downto 0)) * unsigned(b(204 downto 188))); 
temp_mult_45 <= std_logic_vector(unsigned(a(23 downto 0)) * unsigned(b(221 downto 205))); 
temp_mult_46 <= std_logic_vector(unsigned(a(23 downto 0)) * unsigned(b(238 downto 222))); 
temp_mult_47 <= std_logic_vector(unsigned(a(23 downto 0)) * unsigned(b(255 downto 239))); 
temp_mult_48 <= std_logic_vector(unsigned(a(47 downto 24)) * unsigned(b(136 downto 120))); 
temp_mult_49 <= std_logic_vector(unsigned(a(47 downto 24)) * unsigned(b(153 downto 137))); 
temp_mult_50 <= std_logic_vector(unsigned(a(47 downto 24)) * unsigned(b(170 downto 154))); 
temp_mult_51 <= std_logic_vector(unsigned(a(47 downto 24)) * unsigned(b(187 downto 171))); 
temp_mult_52 <= std_logic_vector(unsigned(a(47 downto 24)) * unsigned(b(204 downto 188))); 
temp_mult_53 <= std_logic_vector(unsigned(a(47 downto 24)) * unsigned(b(221 downto 205))); 
temp_mult_54 <= std_logic_vector(unsigned(a(47 downto 24)) * unsigned(b(238 downto 222))); 
temp_mult_55 <= std_logic_vector(unsigned(a(47 downto 24)) * unsigned(b(255 downto 239))); 
temp_mult_56 <= std_logic_vector(unsigned(a(71 downto 48)) * unsigned(b(136 downto 120))); 
temp_mult_57 <= std_logic_vector(unsigned(a(71 downto 48)) * unsigned(b(153 downto 137))); 
temp_mult_58 <= std_logic_vector(unsigned(a(71 downto 48)) * unsigned(b(170 downto 154))); 
temp_mult_59 <= std_logic_vector(unsigned(a(71 downto 48)) * unsigned(b(187 downto 171))); 
temp_mult_60 <= std_logic_vector(unsigned(a(71 downto 48)) * unsigned(b(204 downto 188))); 
temp_mult_61 <= std_logic_vector(unsigned(a(71 downto 48)) * unsigned(b(221 downto 205))); 
temp_mult_62 <= std_logic_vector(unsigned(a(71 downto 48)) * unsigned(b(238 downto 222))); 
temp_mult_63 <= std_logic_vector(unsigned(a(71 downto 48)) * unsigned(b(255 downto 239))); 
temp_mult_64 <= std_logic_vector(unsigned(a(95 downto 72)) * unsigned(b(136 downto 120))); 
temp_mult_65 <= std_logic_vector(unsigned(a(95 downto 72)) * unsigned(b(153 downto 137))); 
temp_mult_66 <= std_logic_vector(unsigned(a(95 downto 72)) * unsigned(b(170 downto 154))); 
temp_mult_67 <= std_logic_vector(unsigned(a(95 downto 72)) * unsigned(b(187 downto 171))); 
temp_mult_68 <= std_logic_vector(unsigned(a(95 downto 72)) * unsigned(b(204 downto 188))); 
temp_mult_69 <= std_logic_vector(unsigned(a(95 downto 72)) * unsigned(b(221 downto 205))); 
temp_mult_70 <= std_logic_vector(unsigned(a(95 downto 72)) * unsigned(b(238 downto 222))); 
temp_mult_71 <= std_logic_vector(unsigned(a(95 downto 72)) * unsigned(b(255 downto 239))); 
temp_mult_72 <= std_logic_vector(unsigned(a(119 downto 96)) * unsigned(b(136 downto 120))); 
temp_mult_73 <= std_logic_vector(unsigned(a(119 downto 96)) * unsigned(b(153 downto 137))); 
temp_mult_74 <= std_logic_vector(unsigned(a(119 downto 96)) * unsigned(b(170 downto 154))); 
temp_mult_75 <= std_logic_vector(unsigned(a(119 downto 96)) * unsigned(b(187 downto 171))); 
temp_mult_76 <= std_logic_vector(unsigned(a(119 downto 96)) * unsigned(b(204 downto 188))); 
temp_mult_77 <= std_logic_vector(unsigned(a(119 downto 96)) * unsigned(b(221 downto 205))); 
temp_mult_78 <= std_logic_vector(unsigned(a(119 downto 96)) * unsigned(b(238 downto 222))); 
temp_mult_79 <= std_logic_vector(unsigned(a(119 downto 96)) * unsigned(b(255 downto 239))); 
temp_mult_80 <= std_logic_vector(unsigned(a(159 downto 136)) * unsigned(b(16 downto 0))); 
temp_mult_81 <= std_logic_vector(unsigned(a(159 downto 136)) * unsigned(b(33 downto 17))); 
temp_mult_82 <= std_logic_vector(unsigned(a(159 downto 136)) * unsigned(b(50 downto 34))); 
temp_mult_83 <= std_logic_vector(unsigned(a(159 downto 136)) * unsigned(b(67 downto 51))); 
temp_mult_84 <= std_logic_vector(unsigned(a(159 downto 136)) * unsigned(b(84 downto 68))); 
temp_mult_85 <= std_logic_vector(unsigned(a(159 downto 136)) * unsigned(b(101 downto 85))); 
temp_mult_86 <= std_logic_vector(unsigned(a(159 downto 136)) * unsigned(b(118 downto 102))); 
temp_mult_87 <= std_logic_vector(unsigned(a(159 downto 136)) * unsigned(b(135 downto 119))); 
temp_mult_88 <= std_logic_vector(unsigned(a(183 downto 160)) * unsigned(b(16 downto 0))); 
temp_mult_89 <= std_logic_vector(unsigned(a(183 downto 160)) * unsigned(b(33 downto 17))); 
temp_mult_90 <= std_logic_vector(unsigned(a(183 downto 160)) * unsigned(b(50 downto 34))); 
temp_mult_91 <= std_logic_vector(unsigned(a(183 downto 160)) * unsigned(b(67 downto 51))); 
temp_mult_92 <= std_logic_vector(unsigned(a(183 downto 160)) * unsigned(b(84 downto 68))); 
temp_mult_93 <= std_logic_vector(unsigned(a(183 downto 160)) * unsigned(b(101 downto 85))); 
temp_mult_94 <= std_logic_vector(unsigned(a(183 downto 160)) * unsigned(b(118 downto 102))); 
temp_mult_95 <= std_logic_vector(unsigned(a(183 downto 160)) * unsigned(b(135 downto 119))); 
temp_mult_96 <= std_logic_vector(unsigned(a(207 downto 184)) * unsigned(b(16 downto 0))); 
temp_mult_97 <= std_logic_vector(unsigned(a(207 downto 184)) * unsigned(b(33 downto 17))); 
temp_mult_98 <= std_logic_vector(unsigned(a(207 downto 184)) * unsigned(b(50 downto 34))); 
temp_mult_99 <= std_logic_vector(unsigned(a(207 downto 184)) * unsigned(b(67 downto 51))); 
temp_mult_100 <= std_logic_vector(unsigned(a(207 downto 184)) * unsigned(b(84 downto 68))); 
temp_mult_101 <= std_logic_vector(unsigned(a(207 downto 184)) * unsigned(b(101 downto 85))); 
temp_mult_102 <= std_logic_vector(unsigned(a(207 downto 184)) * unsigned(b(118 downto 102))); 
temp_mult_103 <= std_logic_vector(unsigned(a(207 downto 184)) * unsigned(b(135 downto 119))); 
temp_mult_104 <= std_logic_vector(unsigned(a(231 downto 208)) * unsigned(b(16 downto 0))); 
temp_mult_105 <= std_logic_vector(unsigned(a(231 downto 208)) * unsigned(b(33 downto 17))); 
temp_mult_106 <= std_logic_vector(unsigned(a(231 downto 208)) * unsigned(b(50 downto 34))); 
temp_mult_107 <= std_logic_vector(unsigned(a(231 downto 208)) * unsigned(b(67 downto 51))); 
temp_mult_108 <= std_logic_vector(unsigned(a(231 downto 208)) * unsigned(b(84 downto 68))); 
temp_mult_109 <= std_logic_vector(unsigned(a(231 downto 208)) * unsigned(b(101 downto 85))); 
temp_mult_110 <= std_logic_vector(unsigned(a(231 downto 208)) * unsigned(b(118 downto 102))); 
temp_mult_111 <= std_logic_vector(unsigned(a(231 downto 208)) * unsigned(b(135 downto 119))); 
temp_mult_112 <= std_logic_vector(unsigned(a(255 downto 232)) * unsigned(b(16 downto 0))); 
temp_mult_113 <= std_logic_vector(unsigned(a(255 downto 232)) * unsigned(b(33 downto 17))); 
temp_mult_114 <= std_logic_vector(unsigned(a(255 downto 232)) * unsigned(b(50 downto 34))); 
temp_mult_115 <= std_logic_vector(unsigned(a(255 downto 232)) * unsigned(b(67 downto 51))); 
temp_mult_116 <= std_logic_vector(unsigned(a(255 downto 232)) * unsigned(b(84 downto 68))); 
temp_mult_117 <= std_logic_vector(unsigned(a(255 downto 232)) * unsigned(b(101 downto 85))); 
temp_mult_118 <= std_logic_vector(unsigned(a(255 downto 232)) * unsigned(b(118 downto 102))); 
temp_mult_119 <= std_logic_vector(unsigned(a(255 downto 232)) * unsigned(b(135 downto 119))); 
temp_mult_120 <= std_logic_vector(unsigned(a(136 downto 120)) * unsigned(b(159 downto 136))); 
temp_mult_121 <= std_logic_vector(unsigned(a(136 downto 120)) * unsigned(b(183 downto 160))); 
temp_mult_122 <= std_logic_vector(unsigned(a(136 downto 120)) * unsigned(b(207 downto 184))); 
temp_mult_123 <= std_logic_vector(unsigned(a(136 downto 120)) * unsigned(b(231 downto 208))); 
temp_mult_124 <= std_logic_vector(unsigned(a(136 downto 120)) * unsigned(b(255 downto 232))); 
temp_mult_125 <= std_logic_vector(unsigned(a(153 downto 137)) * unsigned(b(159 downto 136))); 
temp_mult_126 <= std_logic_vector(unsigned(a(153 downto 137)) * unsigned(b(183 downto 160))); 
temp_mult_127 <= std_logic_vector(unsigned(a(153 downto 137)) * unsigned(b(207 downto 184))); 
temp_mult_128 <= std_logic_vector(unsigned(a(153 downto 137)) * unsigned(b(231 downto 208))); 
temp_mult_129 <= std_logic_vector(unsigned(a(153 downto 137)) * unsigned(b(255 downto 232))); 
temp_mult_130 <= std_logic_vector(unsigned(a(170 downto 154)) * unsigned(b(159 downto 136))); 
temp_mult_131 <= std_logic_vector(unsigned(a(170 downto 154)) * unsigned(b(183 downto 160))); 
temp_mult_132 <= std_logic_vector(unsigned(a(170 downto 154)) * unsigned(b(207 downto 184))); 
temp_mult_133 <= std_logic_vector(unsigned(a(170 downto 154)) * unsigned(b(231 downto 208))); 
temp_mult_134 <= std_logic_vector(unsigned(a(170 downto 154)) * unsigned(b(255 downto 232))); 
temp_mult_135 <= std_logic_vector(unsigned(a(187 downto 171)) * unsigned(b(159 downto 136))); 
temp_mult_136 <= std_logic_vector(unsigned(a(187 downto 171)) * unsigned(b(183 downto 160))); 
temp_mult_137 <= std_logic_vector(unsigned(a(187 downto 171)) * unsigned(b(207 downto 184))); 
temp_mult_138 <= std_logic_vector(unsigned(a(187 downto 171)) * unsigned(b(231 downto 208))); 
temp_mult_139 <= std_logic_vector(unsigned(a(187 downto 171)) * unsigned(b(255 downto 232))); 
temp_mult_140 <= std_logic_vector(unsigned(a(204 downto 188)) * unsigned(b(159 downto 136))); 
temp_mult_141 <= std_logic_vector(unsigned(a(204 downto 188)) * unsigned(b(183 downto 160))); 
temp_mult_142 <= std_logic_vector(unsigned(a(204 downto 188)) * unsigned(b(207 downto 184))); 
temp_mult_143 <= std_logic_vector(unsigned(a(204 downto 188)) * unsigned(b(231 downto 208))); 
temp_mult_144 <= std_logic_vector(unsigned(a(204 downto 188)) * unsigned(b(255 downto 232))); 
temp_mult_145 <= std_logic_vector(unsigned(a(221 downto 205)) * unsigned(b(159 downto 136))); 
temp_mult_146 <= std_logic_vector(unsigned(a(221 downto 205)) * unsigned(b(183 downto 160))); 
temp_mult_147 <= std_logic_vector(unsigned(a(221 downto 205)) * unsigned(b(207 downto 184))); 
temp_mult_148 <= std_logic_vector(unsigned(a(221 downto 205)) * unsigned(b(231 downto 208))); 
temp_mult_149 <= std_logic_vector(unsigned(a(221 downto 205)) * unsigned(b(255 downto 232))); 
temp_mult_150 <= std_logic_vector(unsigned(a(238 downto 222)) * unsigned(b(159 downto 136))); 
temp_mult_151 <= std_logic_vector(unsigned(a(238 downto 222)) * unsigned(b(183 downto 160))); 
temp_mult_152 <= std_logic_vector(unsigned(a(238 downto 222)) * unsigned(b(207 downto 184))); 
temp_mult_153 <= std_logic_vector(unsigned(a(238 downto 222)) * unsigned(b(231 downto 208))); 
temp_mult_154 <= std_logic_vector(unsigned(a(238 downto 222)) * unsigned(b(255 downto 232))); 
temp_mult_155 <= std_logic_vector(unsigned(a(255 downto 239)) * unsigned(b(159 downto 136))); 
temp_mult_156 <= std_logic_vector(unsigned(a(255 downto 239)) * unsigned(b(183 downto 160))); 
temp_mult_157 <= std_logic_vector(unsigned(a(255 downto 239)) * unsigned(b(207 downto 184))); 
temp_mult_158 <= std_logic_vector(unsigned(a(255 downto 239)) * unsigned(b(231 downto 208))); 
temp_mult_159 <= std_logic_vector(unsigned(a(255 downto 239)) * unsigned(b(255 downto 232))); 
temp_mult_160 <= std_logic_vector(unsigned(a(135 downto 120)) * unsigned(b(135 downto 120))); 
temp_part_mult_161 <= (others => a(256));
temp_part_mult_162 <= (others => b(256));
temp_mult_161(511 downto 256) <= temp_part_mult_161 and b(255 downto 0);
temp_mult_161(513 downto 512) <= "00";
temp_mult_162(512 downto 256) <= temp_part_mult_162 and a(256 downto 0); 
temp_mult_162(513) <= temp_mult_162(512); 

partial_product_0(0) <= temp_mult_0(0);
partial_product_0(1) <= temp_mult_0(1);
partial_product_0(2) <= temp_mult_0(2);
partial_product_0(3) <= temp_mult_0(3);
partial_product_0(4) <= temp_mult_0(4);
partial_product_0(5) <= temp_mult_0(5);
partial_product_0(6) <= temp_mult_0(6);
partial_product_0(7) <= temp_mult_0(7);
partial_product_0(8) <= temp_mult_0(8);
partial_product_0(9) <= temp_mult_0(9);
partial_product_0(10) <= temp_mult_0(10);
partial_product_0(11) <= temp_mult_0(11);
partial_product_0(12) <= temp_mult_0(12);
partial_product_0(13) <= temp_mult_0(13);
partial_product_0(14) <= temp_mult_0(14);
partial_product_0(15) <= temp_mult_0(15);
partial_product_0(16) <= temp_mult_0(16);
partial_product_0(17) <= temp_mult_0(17);
partial_product_0(18) <= temp_mult_0(18);
partial_product_0(19) <= temp_mult_0(19);
partial_product_0(20) <= temp_mult_0(20);
partial_product_0(21) <= temp_mult_0(21);
partial_product_0(22) <= temp_mult_0(22);
partial_product_0(23) <= temp_mult_0(23);
partial_product_0(24) <= temp_mult_0(24);
partial_product_0(25) <= temp_mult_0(25);
partial_product_0(26) <= temp_mult_0(26);
partial_product_0(27) <= temp_mult_0(27);
partial_product_0(28) <= temp_mult_0(28);
partial_product_0(29) <= temp_mult_0(29);
partial_product_0(30) <= temp_mult_0(30);
partial_product_0(31) <= temp_mult_0(31);
partial_product_0(32) <= temp_mult_0(32);
partial_product_0(33) <= temp_mult_0(33);
partial_product_0(34) <= temp_mult_0(34);
partial_product_0(35) <= temp_mult_0(35);
partial_product_0(36) <= temp_mult_0(36);
partial_product_0(37) <= temp_mult_0(37);
partial_product_0(38) <= temp_mult_0(38);
partial_product_0(39) <= temp_mult_0(39);
partial_product_0(40) <= temp_mult_0(40);
partial_product_0(41) <= temp_mult_6(41);
partial_product_0(42) <= temp_mult_6(42);
partial_product_0(43) <= temp_mult_6(43);
partial_product_0(44) <= temp_mult_6(44);
partial_product_0(45) <= temp_mult_6(45);
partial_product_0(46) <= temp_mult_6(46);
partial_product_0(47) <= temp_mult_6(47);
partial_product_0(48) <= temp_mult_6(48);
partial_product_0(49) <= temp_mult_6(49);
partial_product_0(50) <= temp_mult_6(50);
partial_product_0(51) <= temp_mult_6(51);
partial_product_0(52) <= temp_mult_6(52);
partial_product_0(53) <= temp_mult_6(53);
partial_product_0(54) <= temp_mult_6(54);
partial_product_0(55) <= temp_mult_6(55);
partial_product_0(56) <= temp_mult_6(56);
partial_product_0(57) <= temp_mult_6(57);
partial_product_0(58) <= temp_mult_6(58);
partial_product_0(59) <= temp_mult_6(59);
partial_product_0(60) <= temp_mult_6(60);
partial_product_0(61) <= temp_mult_6(61);
partial_product_0(62) <= temp_mult_6(62);
partial_product_0(63) <= temp_mult_6(63);
partial_product_0(64) <= temp_mult_6(64);
partial_product_0(65) <= temp_mult_6(65);
partial_product_0(66) <= temp_mult_6(66);
partial_product_0(67) <= temp_mult_6(67);
partial_product_0(68) <= temp_mult_6(68);
partial_product_0(69) <= temp_mult_6(69);
partial_product_0(70) <= temp_mult_6(70);
partial_product_0(71) <= temp_mult_6(71);
partial_product_0(72) <= temp_mult_6(72);
partial_product_0(73) <= temp_mult_6(73);
partial_product_0(74) <= temp_mult_6(74);
partial_product_0(75) <= temp_mult_6(75);
partial_product_0(76) <= temp_mult_6(76);
partial_product_0(77) <= temp_mult_6(77);
partial_product_0(78) <= temp_mult_6(78);
partial_product_0(79) <= temp_mult_6(79);
partial_product_0(80) <= temp_mult_6(80);
partial_product_0(81) <= temp_mult_6(81);
partial_product_0(82) <= temp_mult_12(82);
partial_product_0(83) <= temp_mult_12(83);
partial_product_0(84) <= temp_mult_12(84);
partial_product_0(85) <= temp_mult_12(85);
partial_product_0(86) <= temp_mult_12(86);
partial_product_0(87) <= temp_mult_12(87);
partial_product_0(88) <= temp_mult_12(88);
partial_product_0(89) <= temp_mult_12(89);
partial_product_0(90) <= temp_mult_12(90);
partial_product_0(91) <= temp_mult_12(91);
partial_product_0(92) <= temp_mult_12(92);
partial_product_0(93) <= temp_mult_12(93);
partial_product_0(94) <= temp_mult_12(94);
partial_product_0(95) <= temp_mult_12(95);
partial_product_0(96) <= temp_mult_12(96);
partial_product_0(97) <= temp_mult_12(97);
partial_product_0(98) <= temp_mult_12(98);
partial_product_0(99) <= temp_mult_12(99);
partial_product_0(100) <= temp_mult_12(100);
partial_product_0(101) <= temp_mult_12(101);
partial_product_0(102) <= temp_mult_12(102);
partial_product_0(103) <= temp_mult_12(103);
partial_product_0(104) <= temp_mult_12(104);
partial_product_0(105) <= temp_mult_12(105);
partial_product_0(106) <= temp_mult_12(106);
partial_product_0(107) <= temp_mult_12(107);
partial_product_0(108) <= temp_mult_12(108);
partial_product_0(109) <= temp_mult_12(109);
partial_product_0(110) <= temp_mult_12(110);
partial_product_0(111) <= temp_mult_12(111);
partial_product_0(112) <= temp_mult_12(112);
partial_product_0(113) <= temp_mult_12(113);
partial_product_0(114) <= temp_mult_12(114);
partial_product_0(115) <= temp_mult_12(115);
partial_product_0(116) <= temp_mult_12(116);
partial_product_0(117) <= temp_mult_12(117);
partial_product_0(118) <= temp_mult_12(118);
partial_product_0(119) <= temp_mult_12(119);
partial_product_0(120) <= temp_mult_12(120);
partial_product_0(121) <= temp_mult_12(121);
partial_product_0(122) <= temp_mult_12(122);
partial_product_0(123) <= temp_mult_18(123);
partial_product_0(124) <= temp_mult_18(124);
partial_product_0(125) <= temp_mult_18(125);
partial_product_0(126) <= temp_mult_18(126);
partial_product_0(127) <= temp_mult_18(127);
partial_product_0(128) <= temp_mult_18(128);
partial_product_0(129) <= temp_mult_18(129);
partial_product_0(130) <= temp_mult_18(130);
partial_product_0(131) <= temp_mult_18(131);
partial_product_0(132) <= temp_mult_18(132);
partial_product_0(133) <= temp_mult_18(133);
partial_product_0(134) <= temp_mult_18(134);
partial_product_0(135) <= temp_mult_18(135);
partial_product_0(136) <= temp_mult_18(136);
partial_product_0(137) <= temp_mult_18(137);
partial_product_0(138) <= temp_mult_18(138);
partial_product_0(139) <= temp_mult_18(139);
partial_product_0(140) <= temp_mult_18(140);
partial_product_0(141) <= temp_mult_18(141);
partial_product_0(142) <= temp_mult_18(142);
partial_product_0(143) <= temp_mult_18(143);
partial_product_0(144) <= temp_mult_18(144);
partial_product_0(145) <= temp_mult_18(145);
partial_product_0(146) <= temp_mult_18(146);
partial_product_0(147) <= temp_mult_18(147);
partial_product_0(148) <= temp_mult_18(148);
partial_product_0(149) <= temp_mult_18(149);
partial_product_0(150) <= temp_mult_18(150);
partial_product_0(151) <= temp_mult_18(151);
partial_product_0(152) <= temp_mult_18(152);
partial_product_0(153) <= temp_mult_18(153);
partial_product_0(154) <= temp_mult_18(154);
partial_product_0(155) <= temp_mult_18(155);
partial_product_0(156) <= temp_mult_18(156);
partial_product_0(157) <= temp_mult_18(157);
partial_product_0(158) <= temp_mult_18(158);
partial_product_0(159) <= temp_mult_18(159);
partial_product_0(160) <= temp_mult_18(160);
partial_product_0(161) <= temp_mult_18(161);
partial_product_0(162) <= temp_mult_18(162);
partial_product_0(163) <= temp_mult_18(163);
partial_product_0(164) <= temp_mult_24(164);
partial_product_0(165) <= temp_mult_24(165);
partial_product_0(166) <= temp_mult_24(166);
partial_product_0(167) <= temp_mult_24(167);
partial_product_0(168) <= temp_mult_24(168);
partial_product_0(169) <= temp_mult_24(169);
partial_product_0(170) <= temp_mult_24(170);
partial_product_0(171) <= temp_mult_24(171);
partial_product_0(172) <= temp_mult_24(172);
partial_product_0(173) <= temp_mult_24(173);
partial_product_0(174) <= temp_mult_24(174);
partial_product_0(175) <= temp_mult_24(175);
partial_product_0(176) <= temp_mult_24(176);
partial_product_0(177) <= temp_mult_24(177);
partial_product_0(178) <= temp_mult_24(178);
partial_product_0(179) <= temp_mult_24(179);
partial_product_0(180) <= temp_mult_24(180);
partial_product_0(181) <= temp_mult_24(181);
partial_product_0(182) <= temp_mult_24(182);
partial_product_0(183) <= temp_mult_24(183);
partial_product_0(184) <= temp_mult_24(184);
partial_product_0(185) <= temp_mult_24(185);
partial_product_0(186) <= temp_mult_24(186);
partial_product_0(187) <= temp_mult_24(187);
partial_product_0(188) <= temp_mult_24(188);
partial_product_0(189) <= temp_mult_24(189);
partial_product_0(190) <= temp_mult_24(190);
partial_product_0(191) <= temp_mult_24(191);
partial_product_0(192) <= temp_mult_24(192);
partial_product_0(193) <= temp_mult_24(193);
partial_product_0(194) <= temp_mult_24(194);
partial_product_0(195) <= temp_mult_24(195);
partial_product_0(196) <= temp_mult_24(196);
partial_product_0(197) <= temp_mult_24(197);
partial_product_0(198) <= temp_mult_24(198);
partial_product_0(199) <= temp_mult_24(199);
partial_product_0(200) <= temp_mult_24(200);
partial_product_0(201) <= temp_mult_24(201);
partial_product_0(202) <= temp_mult_24(202);
partial_product_0(203) <= temp_mult_24(203);
partial_product_0(204) <= temp_mult_24(204);
partial_product_0(205) <= temp_mult_45(205);
partial_product_0(206) <= temp_mult_45(206);
partial_product_0(207) <= temp_mult_45(207);
partial_product_0(208) <= temp_mult_45(208);
partial_product_0(209) <= temp_mult_45(209);
partial_product_0(210) <= temp_mult_45(210);
partial_product_0(211) <= temp_mult_45(211);
partial_product_0(212) <= temp_mult_45(212);
partial_product_0(213) <= temp_mult_45(213);
partial_product_0(214) <= temp_mult_45(214);
partial_product_0(215) <= temp_mult_45(215);
partial_product_0(216) <= temp_mult_45(216);
partial_product_0(217) <= temp_mult_45(217);
partial_product_0(218) <= temp_mult_45(218);
partial_product_0(219) <= temp_mult_45(219);
partial_product_0(220) <= temp_mult_45(220);
partial_product_0(221) <= temp_mult_45(221);
partial_product_0(222) <= temp_mult_45(222);
partial_product_0(223) <= temp_mult_45(223);
partial_product_0(224) <= temp_mult_45(224);
partial_product_0(225) <= temp_mult_45(225);
partial_product_0(226) <= temp_mult_45(226);
partial_product_0(227) <= temp_mult_45(227);
partial_product_0(228) <= temp_mult_45(228);
partial_product_0(229) <= temp_mult_45(229);
partial_product_0(230) <= temp_mult_45(230);
partial_product_0(231) <= temp_mult_45(231);
partial_product_0(232) <= temp_mult_45(232);
partial_product_0(233) <= temp_mult_45(233);
partial_product_0(234) <= temp_mult_45(234);
partial_product_0(235) <= temp_mult_45(235);
partial_product_0(236) <= temp_mult_45(236);
partial_product_0(237) <= temp_mult_45(237);
partial_product_0(238) <= temp_mult_45(238);
partial_product_0(239) <= temp_mult_45(239);
partial_product_0(240) <= temp_mult_45(240);
partial_product_0(241) <= temp_mult_45(241);
partial_product_0(242) <= temp_mult_45(242);
partial_product_0(243) <= temp_mult_45(243);
partial_product_0(244) <= temp_mult_45(244);
partial_product_0(245) <= temp_mult_45(245);
partial_product_0(246) <= temp_mult_54(246);
partial_product_0(247) <= temp_mult_54(247);
partial_product_0(248) <= temp_mult_54(248);
partial_product_0(249) <= temp_mult_54(249);
partial_product_0(250) <= temp_mult_54(250);
partial_product_0(251) <= temp_mult_54(251);
partial_product_0(252) <= temp_mult_54(252);
partial_product_0(253) <= temp_mult_54(253);
partial_product_0(254) <= temp_mult_54(254);
partial_product_0(255) <= temp_mult_54(255);
partial_product_0(256) <= temp_mult_54(256);
partial_product_0(257) <= temp_mult_54(257);
partial_product_0(258) <= temp_mult_54(258);
partial_product_0(259) <= temp_mult_54(259);
partial_product_0(260) <= temp_mult_54(260);
partial_product_0(261) <= temp_mult_54(261);
partial_product_0(262) <= temp_mult_54(262);
partial_product_0(263) <= temp_mult_54(263);
partial_product_0(264) <= temp_mult_54(264);
partial_product_0(265) <= temp_mult_54(265);
partial_product_0(266) <= temp_mult_54(266);
partial_product_0(267) <= temp_mult_54(267);
partial_product_0(268) <= temp_mult_54(268);
partial_product_0(269) <= temp_mult_54(269);
partial_product_0(270) <= temp_mult_54(270);
partial_product_0(271) <= temp_mult_54(271);
partial_product_0(272) <= temp_mult_54(272);
partial_product_0(273) <= temp_mult_54(273);
partial_product_0(274) <= temp_mult_54(274);
partial_product_0(275) <= temp_mult_54(275);
partial_product_0(276) <= temp_mult_54(276);
partial_product_0(277) <= temp_mult_54(277);
partial_product_0(278) <= temp_mult_54(278);
partial_product_0(279) <= temp_mult_54(279);
partial_product_0(280) <= temp_mult_54(280);
partial_product_0(281) <= temp_mult_54(281);
partial_product_0(282) <= temp_mult_54(282);
partial_product_0(283) <= temp_mult_54(283);
partial_product_0(284) <= temp_mult_54(284);
partial_product_0(285) <= temp_mult_54(285);
partial_product_0(286) <= temp_mult_54(286);
partial_product_0(287) <= temp_mult_63(287);
partial_product_0(288) <= temp_mult_63(288);
partial_product_0(289) <= temp_mult_63(289);
partial_product_0(290) <= temp_mult_63(290);
partial_product_0(291) <= temp_mult_63(291);
partial_product_0(292) <= temp_mult_63(292);
partial_product_0(293) <= temp_mult_63(293);
partial_product_0(294) <= temp_mult_63(294);
partial_product_0(295) <= temp_mult_63(295);
partial_product_0(296) <= temp_mult_63(296);
partial_product_0(297) <= temp_mult_63(297);
partial_product_0(298) <= temp_mult_63(298);
partial_product_0(299) <= temp_mult_63(299);
partial_product_0(300) <= temp_mult_63(300);
partial_product_0(301) <= temp_mult_63(301);
partial_product_0(302) <= temp_mult_63(302);
partial_product_0(303) <= temp_mult_63(303);
partial_product_0(304) <= temp_mult_63(304);
partial_product_0(305) <= temp_mult_63(305);
partial_product_0(306) <= temp_mult_63(306);
partial_product_0(307) <= temp_mult_63(307);
partial_product_0(308) <= temp_mult_63(308);
partial_product_0(309) <= temp_mult_63(309);
partial_product_0(310) <= temp_mult_63(310);
partial_product_0(311) <= temp_mult_63(311);
partial_product_0(312) <= temp_mult_63(312);
partial_product_0(313) <= temp_mult_63(313);
partial_product_0(314) <= temp_mult_63(314);
partial_product_0(315) <= temp_mult_63(315);
partial_product_0(316) <= temp_mult_63(316);
partial_product_0(317) <= temp_mult_63(317);
partial_product_0(318) <= temp_mult_63(318);
partial_product_0(319) <= temp_mult_63(319);
partial_product_0(320) <= temp_mult_63(320);
partial_product_0(321) <= temp_mult_63(321);
partial_product_0(322) <= temp_mult_63(322);
partial_product_0(323) <= temp_mult_63(323);
partial_product_0(324) <= temp_mult_63(324);
partial_product_0(325) <= temp_mult_63(325);
partial_product_0(326) <= temp_mult_63(326);
partial_product_0(327) <= temp_mult_63(327);
partial_product_0(328) <= temp_mult_123(328);
partial_product_0(329) <= temp_mult_123(329);
partial_product_0(330) <= temp_mult_123(330);
partial_product_0(331) <= temp_mult_123(331);
partial_product_0(332) <= temp_mult_123(332);
partial_product_0(333) <= temp_mult_123(333);
partial_product_0(334) <= temp_mult_123(334);
partial_product_0(335) <= temp_mult_123(335);
partial_product_0(336) <= temp_mult_123(336);
partial_product_0(337) <= temp_mult_123(337);
partial_product_0(338) <= temp_mult_123(338);
partial_product_0(339) <= temp_mult_123(339);
partial_product_0(340) <= temp_mult_123(340);
partial_product_0(341) <= temp_mult_123(341);
partial_product_0(342) <= temp_mult_123(342);
partial_product_0(343) <= temp_mult_123(343);
partial_product_0(344) <= temp_mult_123(344);
partial_product_0(345) <= temp_mult_123(345);
partial_product_0(346) <= temp_mult_123(346);
partial_product_0(347) <= temp_mult_123(347);
partial_product_0(348) <= temp_mult_123(348);
partial_product_0(349) <= temp_mult_123(349);
partial_product_0(350) <= temp_mult_123(350);
partial_product_0(351) <= temp_mult_123(351);
partial_product_0(352) <= temp_mult_123(352);
partial_product_0(353) <= temp_mult_123(353);
partial_product_0(354) <= temp_mult_123(354);
partial_product_0(355) <= temp_mult_123(355);
partial_product_0(356) <= temp_mult_123(356);
partial_product_0(357) <= temp_mult_123(357);
partial_product_0(358) <= temp_mult_123(358);
partial_product_0(359) <= temp_mult_123(359);
partial_product_0(360) <= temp_mult_123(360);
partial_product_0(361) <= temp_mult_123(361);
partial_product_0(362) <= temp_mult_123(362);
partial_product_0(363) <= temp_mult_123(363);
partial_product_0(364) <= temp_mult_123(364);
partial_product_0(365) <= temp_mult_123(365);
partial_product_0(366) <= temp_mult_123(366);
partial_product_0(367) <= temp_mult_123(367);
partial_product_0(368) <= temp_mult_123(368);
partial_product_0(369) <= temp_mult_129(369);
partial_product_0(370) <= temp_mult_129(370);
partial_product_0(371) <= temp_mult_129(371);
partial_product_0(372) <= temp_mult_129(372);
partial_product_0(373) <= temp_mult_129(373);
partial_product_0(374) <= temp_mult_129(374);
partial_product_0(375) <= temp_mult_129(375);
partial_product_0(376) <= temp_mult_129(376);
partial_product_0(377) <= temp_mult_129(377);
partial_product_0(378) <= temp_mult_129(378);
partial_product_0(379) <= temp_mult_129(379);
partial_product_0(380) <= temp_mult_129(380);
partial_product_0(381) <= temp_mult_129(381);
partial_product_0(382) <= temp_mult_129(382);
partial_product_0(383) <= temp_mult_129(383);
partial_product_0(384) <= temp_mult_129(384);
partial_product_0(385) <= temp_mult_129(385);
partial_product_0(386) <= temp_mult_129(386);
partial_product_0(387) <= temp_mult_129(387);
partial_product_0(388) <= temp_mult_129(388);
partial_product_0(389) <= temp_mult_129(389);
partial_product_0(390) <= temp_mult_129(390);
partial_product_0(391) <= temp_mult_129(391);
partial_product_0(392) <= temp_mult_129(392);
partial_product_0(393) <= temp_mult_129(393);
partial_product_0(394) <= temp_mult_129(394);
partial_product_0(395) <= temp_mult_129(395);
partial_product_0(396) <= temp_mult_129(396);
partial_product_0(397) <= temp_mult_129(397);
partial_product_0(398) <= temp_mult_129(398);
partial_product_0(399) <= temp_mult_129(399);
partial_product_0(400) <= temp_mult_129(400);
partial_product_0(401) <= temp_mult_129(401);
partial_product_0(402) <= temp_mult_129(402);
partial_product_0(403) <= temp_mult_129(403);
partial_product_0(404) <= temp_mult_129(404);
partial_product_0(405) <= temp_mult_129(405);
partial_product_0(406) <= temp_mult_129(406);
partial_product_0(407) <= temp_mult_129(407);
partial_product_0(408) <= temp_mult_129(408);
partial_product_0(409) <= temp_mult_129(409);
partial_product_0(410) <= '0';
partial_product_0(411) <= '0';
partial_product_0(412) <= '0';
partial_product_0(413) <= temp_mult_148(413);
partial_product_0(414) <= temp_mult_148(414);
partial_product_0(415) <= temp_mult_148(415);
partial_product_0(416) <= temp_mult_148(416);
partial_product_0(417) <= temp_mult_148(417);
partial_product_0(418) <= temp_mult_148(418);
partial_product_0(419) <= temp_mult_148(419);
partial_product_0(420) <= temp_mult_148(420);
partial_product_0(421) <= temp_mult_148(421);
partial_product_0(422) <= temp_mult_148(422);
partial_product_0(423) <= temp_mult_148(423);
partial_product_0(424) <= temp_mult_148(424);
partial_product_0(425) <= temp_mult_148(425);
partial_product_0(426) <= temp_mult_148(426);
partial_product_0(427) <= temp_mult_148(427);
partial_product_0(428) <= temp_mult_148(428);
partial_product_0(429) <= temp_mult_148(429);
partial_product_0(430) <= temp_mult_148(430);
partial_product_0(431) <= temp_mult_148(431);
partial_product_0(432) <= temp_mult_148(432);
partial_product_0(433) <= temp_mult_148(433);
partial_product_0(434) <= temp_mult_148(434);
partial_product_0(435) <= temp_mult_148(435);
partial_product_0(436) <= temp_mult_148(436);
partial_product_0(437) <= temp_mult_148(437);
partial_product_0(438) <= temp_mult_148(438);
partial_product_0(439) <= temp_mult_148(439);
partial_product_0(440) <= temp_mult_148(440);
partial_product_0(441) <= temp_mult_148(441);
partial_product_0(442) <= temp_mult_148(442);
partial_product_0(443) <= temp_mult_148(443);
partial_product_0(444) <= temp_mult_148(444);
partial_product_0(445) <= temp_mult_148(445);
partial_product_0(446) <= temp_mult_148(446);
partial_product_0(447) <= temp_mult_148(447);
partial_product_0(448) <= temp_mult_148(448);
partial_product_0(449) <= temp_mult_148(449);
partial_product_0(450) <= temp_mult_148(450);
partial_product_0(451) <= temp_mult_148(451);
partial_product_0(452) <= temp_mult_148(452);
partial_product_0(453) <= temp_mult_148(453);
partial_product_0(454) <= temp_mult_154(454);
partial_product_0(455) <= temp_mult_154(455);
partial_product_0(456) <= temp_mult_154(456);
partial_product_0(457) <= temp_mult_154(457);
partial_product_0(458) <= temp_mult_154(458);
partial_product_0(459) <= temp_mult_154(459);
partial_product_0(460) <= temp_mult_154(460);
partial_product_0(461) <= temp_mult_154(461);
partial_product_0(462) <= temp_mult_154(462);
partial_product_0(463) <= temp_mult_154(463);
partial_product_0(464) <= temp_mult_154(464);
partial_product_0(465) <= temp_mult_154(465);
partial_product_0(466) <= temp_mult_154(466);
partial_product_0(467) <= temp_mult_154(467);
partial_product_0(468) <= temp_mult_154(468);
partial_product_0(469) <= temp_mult_154(469);
partial_product_0(470) <= temp_mult_154(470);
partial_product_0(471) <= temp_mult_154(471);
partial_product_0(472) <= temp_mult_154(472);
partial_product_0(473) <= temp_mult_154(473);
partial_product_0(474) <= temp_mult_154(474);
partial_product_0(475) <= temp_mult_154(475);
partial_product_0(476) <= temp_mult_154(476);
partial_product_0(477) <= temp_mult_154(477);
partial_product_0(478) <= temp_mult_154(478);
partial_product_0(479) <= temp_mult_154(479);
partial_product_0(480) <= temp_mult_154(480);
partial_product_0(481) <= temp_mult_154(481);
partial_product_0(482) <= temp_mult_154(482);
partial_product_0(483) <= temp_mult_154(483);
partial_product_0(484) <= temp_mult_154(484);
partial_product_0(485) <= temp_mult_154(485);
partial_product_0(486) <= temp_mult_154(486);
partial_product_0(487) <= temp_mult_154(487);
partial_product_0(488) <= temp_mult_154(488);
partial_product_0(489) <= temp_mult_154(489);
partial_product_0(490) <= temp_mult_154(490);
partial_product_0(491) <= temp_mult_154(491);
partial_product_0(492) <= temp_mult_154(492);
partial_product_0(493) <= temp_mult_154(493);
partial_product_0(494) <= temp_mult_154(494);
partial_product_0(495) <= '0';
partial_product_0(496) <= '0';
partial_product_0(497) <= '0';
partial_product_0(498) <= '0';
partial_product_0(499) <= '0';
partial_product_0(500) <= '0';
partial_product_0(501) <= '0';
partial_product_0(502) <= '0';
partial_product_0(503) <= '0';
partial_product_0(504) <= '0';
partial_product_0(505) <= '0';
partial_product_0(506) <= '0';
partial_product_0(507) <= '0';
partial_product_0(508) <= '0';
partial_product_0(509) <= '0';
partial_product_0(510) <= '0';
partial_product_0(511) <= '0';
partial_product_0(512) <= '0';
partial_product_1(0) <= '0';
partial_product_1(1) <= '0';
partial_product_1(2) <= '0';
partial_product_1(3) <= '0';
partial_product_1(4) <= '0';
partial_product_1(5) <= '0';
partial_product_1(6) <= '0';
partial_product_1(7) <= '0';
partial_product_1(8) <= '0';
partial_product_1(9) <= '0';
partial_product_1(10) <= '0';
partial_product_1(11) <= '0';
partial_product_1(12) <= '0';
partial_product_1(13) <= '0';
partial_product_1(14) <= '0';
partial_product_1(15) <= '0';
partial_product_1(16) <= '0';
partial_product_1(17) <= temp_mult_5(17);
partial_product_1(18) <= temp_mult_5(18);
partial_product_1(19) <= temp_mult_5(19);
partial_product_1(20) <= temp_mult_5(20);
partial_product_1(21) <= temp_mult_5(21);
partial_product_1(22) <= temp_mult_5(22);
partial_product_1(23) <= temp_mult_5(23);
partial_product_1(24) <= temp_mult_5(24);
partial_product_1(25) <= temp_mult_5(25);
partial_product_1(26) <= temp_mult_5(26);
partial_product_1(27) <= temp_mult_5(27);
partial_product_1(28) <= temp_mult_5(28);
partial_product_1(29) <= temp_mult_5(29);
partial_product_1(30) <= temp_mult_5(30);
partial_product_1(31) <= temp_mult_5(31);
partial_product_1(32) <= temp_mult_5(32);
partial_product_1(33) <= temp_mult_5(33);
partial_product_1(34) <= temp_mult_5(34);
partial_product_1(35) <= temp_mult_5(35);
partial_product_1(36) <= temp_mult_5(36);
partial_product_1(37) <= temp_mult_5(37);
partial_product_1(38) <= temp_mult_5(38);
partial_product_1(39) <= temp_mult_5(39);
partial_product_1(40) <= temp_mult_5(40);
partial_product_1(41) <= temp_mult_5(41);
partial_product_1(42) <= temp_mult_5(42);
partial_product_1(43) <= temp_mult_5(43);
partial_product_1(44) <= temp_mult_5(44);
partial_product_1(45) <= temp_mult_5(45);
partial_product_1(46) <= temp_mult_5(46);
partial_product_1(47) <= temp_mult_5(47);
partial_product_1(48) <= temp_mult_5(48);
partial_product_1(49) <= temp_mult_5(49);
partial_product_1(50) <= temp_mult_5(50);
partial_product_1(51) <= temp_mult_5(51);
partial_product_1(52) <= temp_mult_5(52);
partial_product_1(53) <= temp_mult_5(53);
partial_product_1(54) <= temp_mult_5(54);
partial_product_1(55) <= temp_mult_5(55);
partial_product_1(56) <= temp_mult_5(56);
partial_product_1(57) <= temp_mult_5(57);
partial_product_1(58) <= temp_mult_11(58);
partial_product_1(59) <= temp_mult_11(59);
partial_product_1(60) <= temp_mult_11(60);
partial_product_1(61) <= temp_mult_11(61);
partial_product_1(62) <= temp_mult_11(62);
partial_product_1(63) <= temp_mult_11(63);
partial_product_1(64) <= temp_mult_11(64);
partial_product_1(65) <= temp_mult_11(65);
partial_product_1(66) <= temp_mult_11(66);
partial_product_1(67) <= temp_mult_11(67);
partial_product_1(68) <= temp_mult_11(68);
partial_product_1(69) <= temp_mult_11(69);
partial_product_1(70) <= temp_mult_11(70);
partial_product_1(71) <= temp_mult_11(71);
partial_product_1(72) <= temp_mult_11(72);
partial_product_1(73) <= temp_mult_11(73);
partial_product_1(74) <= temp_mult_11(74);
partial_product_1(75) <= temp_mult_11(75);
partial_product_1(76) <= temp_mult_11(76);
partial_product_1(77) <= temp_mult_11(77);
partial_product_1(78) <= temp_mult_11(78);
partial_product_1(79) <= temp_mult_11(79);
partial_product_1(80) <= temp_mult_11(80);
partial_product_1(81) <= temp_mult_11(81);
partial_product_1(82) <= temp_mult_11(82);
partial_product_1(83) <= temp_mult_11(83);
partial_product_1(84) <= temp_mult_11(84);
partial_product_1(85) <= temp_mult_11(85);
partial_product_1(86) <= temp_mult_11(86);
partial_product_1(87) <= temp_mult_11(87);
partial_product_1(88) <= temp_mult_11(88);
partial_product_1(89) <= temp_mult_11(89);
partial_product_1(90) <= temp_mult_11(90);
partial_product_1(91) <= temp_mult_11(91);
partial_product_1(92) <= temp_mult_11(92);
partial_product_1(93) <= temp_mult_11(93);
partial_product_1(94) <= temp_mult_11(94);
partial_product_1(95) <= temp_mult_11(95);
partial_product_1(96) <= temp_mult_11(96);
partial_product_1(97) <= temp_mult_11(97);
partial_product_1(98) <= temp_mult_11(98);
partial_product_1(99) <= temp_mult_17(99);
partial_product_1(100) <= temp_mult_17(100);
partial_product_1(101) <= temp_mult_17(101);
partial_product_1(102) <= temp_mult_17(102);
partial_product_1(103) <= temp_mult_17(103);
partial_product_1(104) <= temp_mult_17(104);
partial_product_1(105) <= temp_mult_17(105);
partial_product_1(106) <= temp_mult_17(106);
partial_product_1(107) <= temp_mult_17(107);
partial_product_1(108) <= temp_mult_17(108);
partial_product_1(109) <= temp_mult_17(109);
partial_product_1(110) <= temp_mult_17(110);
partial_product_1(111) <= temp_mult_17(111);
partial_product_1(112) <= temp_mult_17(112);
partial_product_1(113) <= temp_mult_17(113);
partial_product_1(114) <= temp_mult_17(114);
partial_product_1(115) <= temp_mult_17(115);
partial_product_1(116) <= temp_mult_17(116);
partial_product_1(117) <= temp_mult_17(117);
partial_product_1(118) <= temp_mult_17(118);
partial_product_1(119) <= temp_mult_17(119);
partial_product_1(120) <= temp_mult_17(120);
partial_product_1(121) <= temp_mult_17(121);
partial_product_1(122) <= temp_mult_17(122);
partial_product_1(123) <= temp_mult_17(123);
partial_product_1(124) <= temp_mult_17(124);
partial_product_1(125) <= temp_mult_17(125);
partial_product_1(126) <= temp_mult_17(126);
partial_product_1(127) <= temp_mult_17(127);
partial_product_1(128) <= temp_mult_17(128);
partial_product_1(129) <= temp_mult_17(129);
partial_product_1(130) <= temp_mult_17(130);
partial_product_1(131) <= temp_mult_17(131);
partial_product_1(132) <= temp_mult_17(132);
partial_product_1(133) <= temp_mult_17(133);
partial_product_1(134) <= temp_mult_17(134);
partial_product_1(135) <= temp_mult_17(135);
partial_product_1(136) <= temp_mult_17(136);
partial_product_1(137) <= temp_mult_17(137);
partial_product_1(138) <= temp_mult_17(138);
partial_product_1(139) <= temp_mult_17(139);
partial_product_1(140) <= temp_mult_23(140);
partial_product_1(141) <= temp_mult_23(141);
partial_product_1(142) <= temp_mult_23(142);
partial_product_1(143) <= temp_mult_23(143);
partial_product_1(144) <= temp_mult_23(144);
partial_product_1(145) <= temp_mult_23(145);
partial_product_1(146) <= temp_mult_23(146);
partial_product_1(147) <= temp_mult_23(147);
partial_product_1(148) <= temp_mult_23(148);
partial_product_1(149) <= temp_mult_23(149);
partial_product_1(150) <= temp_mult_23(150);
partial_product_1(151) <= temp_mult_23(151);
partial_product_1(152) <= temp_mult_23(152);
partial_product_1(153) <= temp_mult_23(153);
partial_product_1(154) <= temp_mult_23(154);
partial_product_1(155) <= temp_mult_23(155);
partial_product_1(156) <= temp_mult_23(156);
partial_product_1(157) <= temp_mult_23(157);
partial_product_1(158) <= temp_mult_23(158);
partial_product_1(159) <= temp_mult_23(159);
partial_product_1(160) <= temp_mult_23(160);
partial_product_1(161) <= temp_mult_23(161);
partial_product_1(162) <= temp_mult_23(162);
partial_product_1(163) <= temp_mult_23(163);
partial_product_1(164) <= temp_mult_23(164);
partial_product_1(165) <= temp_mult_23(165);
partial_product_1(166) <= temp_mult_23(166);
partial_product_1(167) <= temp_mult_23(167);
partial_product_1(168) <= temp_mult_23(168);
partial_product_1(169) <= temp_mult_23(169);
partial_product_1(170) <= temp_mult_23(170);
partial_product_1(171) <= temp_mult_23(171);
partial_product_1(172) <= temp_mult_23(172);
partial_product_1(173) <= temp_mult_23(173);
partial_product_1(174) <= temp_mult_23(174);
partial_product_1(175) <= temp_mult_23(175);
partial_product_1(176) <= temp_mult_23(176);
partial_product_1(177) <= temp_mult_23(177);
partial_product_1(178) <= temp_mult_23(178);
partial_product_1(179) <= temp_mult_23(179);
partial_product_1(180) <= temp_mult_23(180);
partial_product_1(181) <= temp_mult_29(181);
partial_product_1(182) <= temp_mult_29(182);
partial_product_1(183) <= temp_mult_29(183);
partial_product_1(184) <= temp_mult_29(184);
partial_product_1(185) <= temp_mult_29(185);
partial_product_1(186) <= temp_mult_29(186);
partial_product_1(187) <= temp_mult_29(187);
partial_product_1(188) <= temp_mult_29(188);
partial_product_1(189) <= temp_mult_29(189);
partial_product_1(190) <= temp_mult_29(190);
partial_product_1(191) <= temp_mult_29(191);
partial_product_1(192) <= temp_mult_29(192);
partial_product_1(193) <= temp_mult_29(193);
partial_product_1(194) <= temp_mult_29(194);
partial_product_1(195) <= temp_mult_29(195);
partial_product_1(196) <= temp_mult_29(196);
partial_product_1(197) <= temp_mult_29(197);
partial_product_1(198) <= temp_mult_29(198);
partial_product_1(199) <= temp_mult_29(199);
partial_product_1(200) <= temp_mult_29(200);
partial_product_1(201) <= temp_mult_29(201);
partial_product_1(202) <= temp_mult_29(202);
partial_product_1(203) <= temp_mult_29(203);
partial_product_1(204) <= temp_mult_29(204);
partial_product_1(205) <= temp_mult_29(205);
partial_product_1(206) <= temp_mult_29(206);
partial_product_1(207) <= temp_mult_29(207);
partial_product_1(208) <= temp_mult_29(208);
partial_product_1(209) <= temp_mult_29(209);
partial_product_1(210) <= temp_mult_29(210);
partial_product_1(211) <= temp_mult_29(211);
partial_product_1(212) <= temp_mult_29(212);
partial_product_1(213) <= temp_mult_29(213);
partial_product_1(214) <= temp_mult_29(214);
partial_product_1(215) <= temp_mult_29(215);
partial_product_1(216) <= temp_mult_29(216);
partial_product_1(217) <= temp_mult_29(217);
partial_product_1(218) <= temp_mult_29(218);
partial_product_1(219) <= temp_mult_29(219);
partial_product_1(220) <= temp_mult_29(220);
partial_product_1(221) <= temp_mult_29(221);
partial_product_1(222) <= temp_mult_46(222);
partial_product_1(223) <= temp_mult_46(223);
partial_product_1(224) <= temp_mult_46(224);
partial_product_1(225) <= temp_mult_46(225);
partial_product_1(226) <= temp_mult_46(226);
partial_product_1(227) <= temp_mult_46(227);
partial_product_1(228) <= temp_mult_46(228);
partial_product_1(229) <= temp_mult_46(229);
partial_product_1(230) <= temp_mult_46(230);
partial_product_1(231) <= temp_mult_46(231);
partial_product_1(232) <= temp_mult_46(232);
partial_product_1(233) <= temp_mult_46(233);
partial_product_1(234) <= temp_mult_46(234);
partial_product_1(235) <= temp_mult_46(235);
partial_product_1(236) <= temp_mult_46(236);
partial_product_1(237) <= temp_mult_46(237);
partial_product_1(238) <= temp_mult_46(238);
partial_product_1(239) <= temp_mult_46(239);
partial_product_1(240) <= temp_mult_46(240);
partial_product_1(241) <= temp_mult_46(241);
partial_product_1(242) <= temp_mult_46(242);
partial_product_1(243) <= temp_mult_46(243);
partial_product_1(244) <= temp_mult_46(244);
partial_product_1(245) <= temp_mult_46(245);
partial_product_1(246) <= temp_mult_46(246);
partial_product_1(247) <= temp_mult_46(247);
partial_product_1(248) <= temp_mult_46(248);
partial_product_1(249) <= temp_mult_46(249);
partial_product_1(250) <= temp_mult_46(250);
partial_product_1(251) <= temp_mult_46(251);
partial_product_1(252) <= temp_mult_46(252);
partial_product_1(253) <= temp_mult_46(253);
partial_product_1(254) <= temp_mult_46(254);
partial_product_1(255) <= temp_mult_46(255);
partial_product_1(256) <= temp_mult_46(256);
partial_product_1(257) <= temp_mult_46(257);
partial_product_1(258) <= temp_mult_46(258);
partial_product_1(259) <= temp_mult_46(259);
partial_product_1(260) <= temp_mult_46(260);
partial_product_1(261) <= temp_mult_46(261);
partial_product_1(262) <= temp_mult_46(262);
partial_product_1(263) <= temp_mult_55(263);
partial_product_1(264) <= temp_mult_55(264);
partial_product_1(265) <= temp_mult_55(265);
partial_product_1(266) <= temp_mult_55(266);
partial_product_1(267) <= temp_mult_55(267);
partial_product_1(268) <= temp_mult_55(268);
partial_product_1(269) <= temp_mult_55(269);
partial_product_1(270) <= temp_mult_55(270);
partial_product_1(271) <= temp_mult_55(271);
partial_product_1(272) <= temp_mult_55(272);
partial_product_1(273) <= temp_mult_55(273);
partial_product_1(274) <= temp_mult_55(274);
partial_product_1(275) <= temp_mult_55(275);
partial_product_1(276) <= temp_mult_55(276);
partial_product_1(277) <= temp_mult_55(277);
partial_product_1(278) <= temp_mult_55(278);
partial_product_1(279) <= temp_mult_55(279);
partial_product_1(280) <= temp_mult_55(280);
partial_product_1(281) <= temp_mult_55(281);
partial_product_1(282) <= temp_mult_55(282);
partial_product_1(283) <= temp_mult_55(283);
partial_product_1(284) <= temp_mult_55(284);
partial_product_1(285) <= temp_mult_55(285);
partial_product_1(286) <= temp_mult_55(286);
partial_product_1(287) <= temp_mult_55(287);
partial_product_1(288) <= temp_mult_55(288);
partial_product_1(289) <= temp_mult_55(289);
partial_product_1(290) <= temp_mult_55(290);
partial_product_1(291) <= temp_mult_55(291);
partial_product_1(292) <= temp_mult_55(292);
partial_product_1(293) <= temp_mult_55(293);
partial_product_1(294) <= temp_mult_55(294);
partial_product_1(295) <= temp_mult_55(295);
partial_product_1(296) <= temp_mult_55(296);
partial_product_1(297) <= temp_mult_55(297);
partial_product_1(298) <= temp_mult_55(298);
partial_product_1(299) <= temp_mult_55(299);
partial_product_1(300) <= temp_mult_55(300);
partial_product_1(301) <= temp_mult_55(301);
partial_product_1(302) <= temp_mult_55(302);
partial_product_1(303) <= temp_mult_55(303);
partial_product_1(304) <= temp_mult_122(304);
partial_product_1(305) <= temp_mult_122(305);
partial_product_1(306) <= temp_mult_122(306);
partial_product_1(307) <= temp_mult_122(307);
partial_product_1(308) <= temp_mult_122(308);
partial_product_1(309) <= temp_mult_122(309);
partial_product_1(310) <= temp_mult_122(310);
partial_product_1(311) <= temp_mult_122(311);
partial_product_1(312) <= temp_mult_122(312);
partial_product_1(313) <= temp_mult_122(313);
partial_product_1(314) <= temp_mult_122(314);
partial_product_1(315) <= temp_mult_122(315);
partial_product_1(316) <= temp_mult_122(316);
partial_product_1(317) <= temp_mult_122(317);
partial_product_1(318) <= temp_mult_122(318);
partial_product_1(319) <= temp_mult_122(319);
partial_product_1(320) <= temp_mult_122(320);
partial_product_1(321) <= temp_mult_122(321);
partial_product_1(322) <= temp_mult_122(322);
partial_product_1(323) <= temp_mult_122(323);
partial_product_1(324) <= temp_mult_122(324);
partial_product_1(325) <= temp_mult_122(325);
partial_product_1(326) <= temp_mult_122(326);
partial_product_1(327) <= temp_mult_122(327);
partial_product_1(328) <= temp_mult_122(328);
partial_product_1(329) <= temp_mult_122(329);
partial_product_1(330) <= temp_mult_122(330);
partial_product_1(331) <= temp_mult_122(331);
partial_product_1(332) <= temp_mult_122(332);
partial_product_1(333) <= temp_mult_122(333);
partial_product_1(334) <= temp_mult_122(334);
partial_product_1(335) <= temp_mult_122(335);
partial_product_1(336) <= temp_mult_122(336);
partial_product_1(337) <= temp_mult_122(337);
partial_product_1(338) <= temp_mult_122(338);
partial_product_1(339) <= temp_mult_122(339);
partial_product_1(340) <= temp_mult_122(340);
partial_product_1(341) <= temp_mult_122(341);
partial_product_1(342) <= temp_mult_122(342);
partial_product_1(343) <= temp_mult_122(343);
partial_product_1(344) <= temp_mult_122(344);
partial_product_1(345) <= temp_mult_128(345);
partial_product_1(346) <= temp_mult_128(346);
partial_product_1(347) <= temp_mult_128(347);
partial_product_1(348) <= temp_mult_128(348);
partial_product_1(349) <= temp_mult_128(349);
partial_product_1(350) <= temp_mult_128(350);
partial_product_1(351) <= temp_mult_128(351);
partial_product_1(352) <= temp_mult_128(352);
partial_product_1(353) <= temp_mult_128(353);
partial_product_1(354) <= temp_mult_128(354);
partial_product_1(355) <= temp_mult_128(355);
partial_product_1(356) <= temp_mult_128(356);
partial_product_1(357) <= temp_mult_128(357);
partial_product_1(358) <= temp_mult_128(358);
partial_product_1(359) <= temp_mult_128(359);
partial_product_1(360) <= temp_mult_128(360);
partial_product_1(361) <= temp_mult_128(361);
partial_product_1(362) <= temp_mult_128(362);
partial_product_1(363) <= temp_mult_128(363);
partial_product_1(364) <= temp_mult_128(364);
partial_product_1(365) <= temp_mult_128(365);
partial_product_1(366) <= temp_mult_128(366);
partial_product_1(367) <= temp_mult_128(367);
partial_product_1(368) <= temp_mult_128(368);
partial_product_1(369) <= temp_mult_128(369);
partial_product_1(370) <= temp_mult_128(370);
partial_product_1(371) <= temp_mult_128(371);
partial_product_1(372) <= temp_mult_128(372);
partial_product_1(373) <= temp_mult_128(373);
partial_product_1(374) <= temp_mult_128(374);
partial_product_1(375) <= temp_mult_128(375);
partial_product_1(376) <= temp_mult_128(376);
partial_product_1(377) <= temp_mult_128(377);
partial_product_1(378) <= temp_mult_128(378);
partial_product_1(379) <= temp_mult_128(379);
partial_product_1(380) <= temp_mult_128(380);
partial_product_1(381) <= temp_mult_128(381);
partial_product_1(382) <= temp_mult_128(382);
partial_product_1(383) <= temp_mult_128(383);
partial_product_1(384) <= temp_mult_128(384);
partial_product_1(385) <= temp_mult_128(385);
partial_product_1(386) <= temp_mult_134(386);
partial_product_1(387) <= temp_mult_134(387);
partial_product_1(388) <= temp_mult_134(388);
partial_product_1(389) <= temp_mult_134(389);
partial_product_1(390) <= temp_mult_134(390);
partial_product_1(391) <= temp_mult_134(391);
partial_product_1(392) <= temp_mult_134(392);
partial_product_1(393) <= temp_mult_134(393);
partial_product_1(394) <= temp_mult_134(394);
partial_product_1(395) <= temp_mult_134(395);
partial_product_1(396) <= temp_mult_134(396);
partial_product_1(397) <= temp_mult_134(397);
partial_product_1(398) <= temp_mult_134(398);
partial_product_1(399) <= temp_mult_134(399);
partial_product_1(400) <= temp_mult_134(400);
partial_product_1(401) <= temp_mult_134(401);
partial_product_1(402) <= temp_mult_134(402);
partial_product_1(403) <= temp_mult_134(403);
partial_product_1(404) <= temp_mult_134(404);
partial_product_1(405) <= temp_mult_134(405);
partial_product_1(406) <= temp_mult_134(406);
partial_product_1(407) <= temp_mult_134(407);
partial_product_1(408) <= temp_mult_134(408);
partial_product_1(409) <= temp_mult_134(409);
partial_product_1(410) <= temp_mult_134(410);
partial_product_1(411) <= temp_mult_134(411);
partial_product_1(412) <= temp_mult_134(412);
partial_product_1(413) <= temp_mult_134(413);
partial_product_1(414) <= temp_mult_134(414);
partial_product_1(415) <= temp_mult_134(415);
partial_product_1(416) <= temp_mult_134(416);
partial_product_1(417) <= temp_mult_134(417);
partial_product_1(418) <= temp_mult_134(418);
partial_product_1(419) <= temp_mult_134(419);
partial_product_1(420) <= temp_mult_134(420);
partial_product_1(421) <= temp_mult_134(421);
partial_product_1(422) <= temp_mult_134(422);
partial_product_1(423) <= temp_mult_134(423);
partial_product_1(424) <= temp_mult_134(424);
partial_product_1(425) <= temp_mult_134(425);
partial_product_1(426) <= temp_mult_134(426);
partial_product_1(427) <= '0';
partial_product_1(428) <= '0';
partial_product_1(429) <= '0';
partial_product_1(430) <= temp_mult_153(430);
partial_product_1(431) <= temp_mult_153(431);
partial_product_1(432) <= temp_mult_153(432);
partial_product_1(433) <= temp_mult_153(433);
partial_product_1(434) <= temp_mult_153(434);
partial_product_1(435) <= temp_mult_153(435);
partial_product_1(436) <= temp_mult_153(436);
partial_product_1(437) <= temp_mult_153(437);
partial_product_1(438) <= temp_mult_153(438);
partial_product_1(439) <= temp_mult_153(439);
partial_product_1(440) <= temp_mult_153(440);
partial_product_1(441) <= temp_mult_153(441);
partial_product_1(442) <= temp_mult_153(442);
partial_product_1(443) <= temp_mult_153(443);
partial_product_1(444) <= temp_mult_153(444);
partial_product_1(445) <= temp_mult_153(445);
partial_product_1(446) <= temp_mult_153(446);
partial_product_1(447) <= temp_mult_153(447);
partial_product_1(448) <= temp_mult_153(448);
partial_product_1(449) <= temp_mult_153(449);
partial_product_1(450) <= temp_mult_153(450);
partial_product_1(451) <= temp_mult_153(451);
partial_product_1(452) <= temp_mult_153(452);
partial_product_1(453) <= temp_mult_153(453);
partial_product_1(454) <= temp_mult_153(454);
partial_product_1(455) <= temp_mult_153(455);
partial_product_1(456) <= temp_mult_153(456);
partial_product_1(457) <= temp_mult_153(457);
partial_product_1(458) <= temp_mult_153(458);
partial_product_1(459) <= temp_mult_153(459);
partial_product_1(460) <= temp_mult_153(460);
partial_product_1(461) <= temp_mult_153(461);
partial_product_1(462) <= temp_mult_153(462);
partial_product_1(463) <= temp_mult_153(463);
partial_product_1(464) <= temp_mult_153(464);
partial_product_1(465) <= temp_mult_153(465);
partial_product_1(466) <= temp_mult_153(466);
partial_product_1(467) <= temp_mult_153(467);
partial_product_1(468) <= temp_mult_153(468);
partial_product_1(469) <= temp_mult_153(469);
partial_product_1(470) <= temp_mult_153(470);
partial_product_1(471) <= temp_mult_159(471);
partial_product_1(472) <= temp_mult_159(472);
partial_product_1(473) <= temp_mult_159(473);
partial_product_1(474) <= temp_mult_159(474);
partial_product_1(475) <= temp_mult_159(475);
partial_product_1(476) <= temp_mult_159(476);
partial_product_1(477) <= temp_mult_159(477);
partial_product_1(478) <= temp_mult_159(478);
partial_product_1(479) <= temp_mult_159(479);
partial_product_1(480) <= temp_mult_159(480);
partial_product_1(481) <= temp_mult_159(481);
partial_product_1(482) <= temp_mult_159(482);
partial_product_1(483) <= temp_mult_159(483);
partial_product_1(484) <= temp_mult_159(484);
partial_product_1(485) <= temp_mult_159(485);
partial_product_1(486) <= temp_mult_159(486);
partial_product_1(487) <= temp_mult_159(487);
partial_product_1(488) <= temp_mult_159(488);
partial_product_1(489) <= temp_mult_159(489);
partial_product_1(490) <= temp_mult_159(490);
partial_product_1(491) <= temp_mult_159(491);
partial_product_1(492) <= temp_mult_159(492);
partial_product_1(493) <= temp_mult_159(493);
partial_product_1(494) <= temp_mult_159(494);
partial_product_1(495) <= temp_mult_159(495);
partial_product_1(496) <= temp_mult_159(496);
partial_product_1(497) <= temp_mult_159(497);
partial_product_1(498) <= temp_mult_159(498);
partial_product_1(499) <= temp_mult_159(499);
partial_product_1(500) <= temp_mult_159(500);
partial_product_1(501) <= temp_mult_159(501);
partial_product_1(502) <= temp_mult_159(502);
partial_product_1(503) <= temp_mult_159(503);
partial_product_1(504) <= temp_mult_159(504);
partial_product_1(505) <= temp_mult_159(505);
partial_product_1(506) <= temp_mult_159(506);
partial_product_1(507) <= temp_mult_159(507);
partial_product_1(508) <= temp_mult_159(508);
partial_product_1(509) <= temp_mult_159(509);
partial_product_1(510) <= temp_mult_159(510);
partial_product_1(511) <= temp_mult_159(511);
partial_product_1(512) <= '0';
partial_product_2(0) <= '0';
partial_product_2(1) <= '0';
partial_product_2(2) <= '0';
partial_product_2(3) <= '0';
partial_product_2(4) <= '0';
partial_product_2(5) <= '0';
partial_product_2(6) <= '0';
partial_product_2(7) <= '0';
partial_product_2(8) <= '0';
partial_product_2(9) <= '0';
partial_product_2(10) <= '0';
partial_product_2(11) <= '0';
partial_product_2(12) <= '0';
partial_product_2(13) <= '0';
partial_product_2(14) <= '0';
partial_product_2(15) <= '0';
partial_product_2(16) <= '0';
partial_product_2(17) <= '0';
partial_product_2(18) <= '0';
partial_product_2(19) <= '0';
partial_product_2(20) <= '0';
partial_product_2(21) <= '0';
partial_product_2(22) <= '0';
partial_product_2(23) <= '0';
partial_product_2(24) <= temp_mult_1(24);
partial_product_2(25) <= temp_mult_1(25);
partial_product_2(26) <= temp_mult_1(26);
partial_product_2(27) <= temp_mult_1(27);
partial_product_2(28) <= temp_mult_1(28);
partial_product_2(29) <= temp_mult_1(29);
partial_product_2(30) <= temp_mult_1(30);
partial_product_2(31) <= temp_mult_1(31);
partial_product_2(32) <= temp_mult_1(32);
partial_product_2(33) <= temp_mult_1(33);
partial_product_2(34) <= temp_mult_1(34);
partial_product_2(35) <= temp_mult_1(35);
partial_product_2(36) <= temp_mult_1(36);
partial_product_2(37) <= temp_mult_1(37);
partial_product_2(38) <= temp_mult_1(38);
partial_product_2(39) <= temp_mult_1(39);
partial_product_2(40) <= temp_mult_1(40);
partial_product_2(41) <= temp_mult_1(41);
partial_product_2(42) <= temp_mult_1(42);
partial_product_2(43) <= temp_mult_1(43);
partial_product_2(44) <= temp_mult_1(44);
partial_product_2(45) <= temp_mult_1(45);
partial_product_2(46) <= temp_mult_1(46);
partial_product_2(47) <= temp_mult_1(47);
partial_product_2(48) <= temp_mult_1(48);
partial_product_2(49) <= temp_mult_1(49);
partial_product_2(50) <= temp_mult_1(50);
partial_product_2(51) <= temp_mult_1(51);
partial_product_2(52) <= temp_mult_1(52);
partial_product_2(53) <= temp_mult_1(53);
partial_product_2(54) <= temp_mult_1(54);
partial_product_2(55) <= temp_mult_1(55);
partial_product_2(56) <= temp_mult_1(56);
partial_product_2(57) <= temp_mult_1(57);
partial_product_2(58) <= temp_mult_1(58);
partial_product_2(59) <= temp_mult_1(59);
partial_product_2(60) <= temp_mult_1(60);
partial_product_2(61) <= temp_mult_1(61);
partial_product_2(62) <= temp_mult_1(62);
partial_product_2(63) <= temp_mult_1(63);
partial_product_2(64) <= temp_mult_1(64);
partial_product_2(65) <= temp_mult_7(65);
partial_product_2(66) <= temp_mult_7(66);
partial_product_2(67) <= temp_mult_7(67);
partial_product_2(68) <= temp_mult_7(68);
partial_product_2(69) <= temp_mult_7(69);
partial_product_2(70) <= temp_mult_7(70);
partial_product_2(71) <= temp_mult_7(71);
partial_product_2(72) <= temp_mult_7(72);
partial_product_2(73) <= temp_mult_7(73);
partial_product_2(74) <= temp_mult_7(74);
partial_product_2(75) <= temp_mult_7(75);
partial_product_2(76) <= temp_mult_7(76);
partial_product_2(77) <= temp_mult_7(77);
partial_product_2(78) <= temp_mult_7(78);
partial_product_2(79) <= temp_mult_7(79);
partial_product_2(80) <= temp_mult_7(80);
partial_product_2(81) <= temp_mult_7(81);
partial_product_2(82) <= temp_mult_7(82);
partial_product_2(83) <= temp_mult_7(83);
partial_product_2(84) <= temp_mult_7(84);
partial_product_2(85) <= temp_mult_7(85);
partial_product_2(86) <= temp_mult_7(86);
partial_product_2(87) <= temp_mult_7(87);
partial_product_2(88) <= temp_mult_7(88);
partial_product_2(89) <= temp_mult_7(89);
partial_product_2(90) <= temp_mult_7(90);
partial_product_2(91) <= temp_mult_7(91);
partial_product_2(92) <= temp_mult_7(92);
partial_product_2(93) <= temp_mult_7(93);
partial_product_2(94) <= temp_mult_7(94);
partial_product_2(95) <= temp_mult_7(95);
partial_product_2(96) <= temp_mult_7(96);
partial_product_2(97) <= temp_mult_7(97);
partial_product_2(98) <= temp_mult_7(98);
partial_product_2(99) <= temp_mult_7(99);
partial_product_2(100) <= temp_mult_7(100);
partial_product_2(101) <= temp_mult_7(101);
partial_product_2(102) <= temp_mult_7(102);
partial_product_2(103) <= temp_mult_7(103);
partial_product_2(104) <= temp_mult_7(104);
partial_product_2(105) <= temp_mult_7(105);
partial_product_2(106) <= temp_mult_13(106);
partial_product_2(107) <= temp_mult_13(107);
partial_product_2(108) <= temp_mult_13(108);
partial_product_2(109) <= temp_mult_13(109);
partial_product_2(110) <= temp_mult_13(110);
partial_product_2(111) <= temp_mult_13(111);
partial_product_2(112) <= temp_mult_13(112);
partial_product_2(113) <= temp_mult_13(113);
partial_product_2(114) <= temp_mult_13(114);
partial_product_2(115) <= temp_mult_13(115);
partial_product_2(116) <= temp_mult_13(116);
partial_product_2(117) <= temp_mult_13(117);
partial_product_2(118) <= temp_mult_13(118);
partial_product_2(119) <= temp_mult_13(119);
partial_product_2(120) <= temp_mult_13(120);
partial_product_2(121) <= temp_mult_13(121);
partial_product_2(122) <= temp_mult_13(122);
partial_product_2(123) <= temp_mult_13(123);
partial_product_2(124) <= temp_mult_13(124);
partial_product_2(125) <= temp_mult_13(125);
partial_product_2(126) <= temp_mult_13(126);
partial_product_2(127) <= temp_mult_13(127);
partial_product_2(128) <= temp_mult_13(128);
partial_product_2(129) <= temp_mult_13(129);
partial_product_2(130) <= temp_mult_13(130);
partial_product_2(131) <= temp_mult_13(131);
partial_product_2(132) <= temp_mult_13(132);
partial_product_2(133) <= temp_mult_13(133);
partial_product_2(134) <= temp_mult_13(134);
partial_product_2(135) <= temp_mult_13(135);
partial_product_2(136) <= temp_mult_13(136);
partial_product_2(137) <= temp_mult_13(137);
partial_product_2(138) <= temp_mult_13(138);
partial_product_2(139) <= temp_mult_13(139);
partial_product_2(140) <= temp_mult_13(140);
partial_product_2(141) <= temp_mult_13(141);
partial_product_2(142) <= temp_mult_13(142);
partial_product_2(143) <= temp_mult_13(143);
partial_product_2(144) <= temp_mult_13(144);
partial_product_2(145) <= temp_mult_13(145);
partial_product_2(146) <= temp_mult_13(146);
partial_product_2(147) <= temp_mult_19(147);
partial_product_2(148) <= temp_mult_19(148);
partial_product_2(149) <= temp_mult_19(149);
partial_product_2(150) <= temp_mult_19(150);
partial_product_2(151) <= temp_mult_19(151);
partial_product_2(152) <= temp_mult_19(152);
partial_product_2(153) <= temp_mult_19(153);
partial_product_2(154) <= temp_mult_19(154);
partial_product_2(155) <= temp_mult_19(155);
partial_product_2(156) <= temp_mult_19(156);
partial_product_2(157) <= temp_mult_19(157);
partial_product_2(158) <= temp_mult_19(158);
partial_product_2(159) <= temp_mult_19(159);
partial_product_2(160) <= temp_mult_19(160);
partial_product_2(161) <= temp_mult_19(161);
partial_product_2(162) <= temp_mult_19(162);
partial_product_2(163) <= temp_mult_19(163);
partial_product_2(164) <= temp_mult_19(164);
partial_product_2(165) <= temp_mult_19(165);
partial_product_2(166) <= temp_mult_19(166);
partial_product_2(167) <= temp_mult_19(167);
partial_product_2(168) <= temp_mult_19(168);
partial_product_2(169) <= temp_mult_19(169);
partial_product_2(170) <= temp_mult_19(170);
partial_product_2(171) <= temp_mult_19(171);
partial_product_2(172) <= temp_mult_19(172);
partial_product_2(173) <= temp_mult_19(173);
partial_product_2(174) <= temp_mult_19(174);
partial_product_2(175) <= temp_mult_19(175);
partial_product_2(176) <= temp_mult_19(176);
partial_product_2(177) <= temp_mult_19(177);
partial_product_2(178) <= temp_mult_19(178);
partial_product_2(179) <= temp_mult_19(179);
partial_product_2(180) <= temp_mult_19(180);
partial_product_2(181) <= temp_mult_19(181);
partial_product_2(182) <= temp_mult_19(182);
partial_product_2(183) <= temp_mult_19(183);
partial_product_2(184) <= temp_mult_19(184);
partial_product_2(185) <= temp_mult_19(185);
partial_product_2(186) <= temp_mult_19(186);
partial_product_2(187) <= temp_mult_19(187);
partial_product_2(188) <= temp_mult_44(188);
partial_product_2(189) <= temp_mult_44(189);
partial_product_2(190) <= temp_mult_44(190);
partial_product_2(191) <= temp_mult_44(191);
partial_product_2(192) <= temp_mult_44(192);
partial_product_2(193) <= temp_mult_44(193);
partial_product_2(194) <= temp_mult_44(194);
partial_product_2(195) <= temp_mult_44(195);
partial_product_2(196) <= temp_mult_44(196);
partial_product_2(197) <= temp_mult_44(197);
partial_product_2(198) <= temp_mult_44(198);
partial_product_2(199) <= temp_mult_44(199);
partial_product_2(200) <= temp_mult_44(200);
partial_product_2(201) <= temp_mult_44(201);
partial_product_2(202) <= temp_mult_44(202);
partial_product_2(203) <= temp_mult_44(203);
partial_product_2(204) <= temp_mult_44(204);
partial_product_2(205) <= temp_mult_44(205);
partial_product_2(206) <= temp_mult_44(206);
partial_product_2(207) <= temp_mult_44(207);
partial_product_2(208) <= temp_mult_44(208);
partial_product_2(209) <= temp_mult_44(209);
partial_product_2(210) <= temp_mult_44(210);
partial_product_2(211) <= temp_mult_44(211);
partial_product_2(212) <= temp_mult_44(212);
partial_product_2(213) <= temp_mult_44(213);
partial_product_2(214) <= temp_mult_44(214);
partial_product_2(215) <= temp_mult_44(215);
partial_product_2(216) <= temp_mult_44(216);
partial_product_2(217) <= temp_mult_44(217);
partial_product_2(218) <= temp_mult_44(218);
partial_product_2(219) <= temp_mult_44(219);
partial_product_2(220) <= temp_mult_44(220);
partial_product_2(221) <= temp_mult_44(221);
partial_product_2(222) <= temp_mult_44(222);
partial_product_2(223) <= temp_mult_44(223);
partial_product_2(224) <= temp_mult_44(224);
partial_product_2(225) <= temp_mult_44(225);
partial_product_2(226) <= temp_mult_44(226);
partial_product_2(227) <= temp_mult_44(227);
partial_product_2(228) <= temp_mult_44(228);
partial_product_2(229) <= temp_mult_53(229);
partial_product_2(230) <= temp_mult_53(230);
partial_product_2(231) <= temp_mult_53(231);
partial_product_2(232) <= temp_mult_53(232);
partial_product_2(233) <= temp_mult_53(233);
partial_product_2(234) <= temp_mult_53(234);
partial_product_2(235) <= temp_mult_53(235);
partial_product_2(236) <= temp_mult_53(236);
partial_product_2(237) <= temp_mult_53(237);
partial_product_2(238) <= temp_mult_53(238);
partial_product_2(239) <= temp_mult_53(239);
partial_product_2(240) <= temp_mult_53(240);
partial_product_2(241) <= temp_mult_53(241);
partial_product_2(242) <= temp_mult_53(242);
partial_product_2(243) <= temp_mult_53(243);
partial_product_2(244) <= temp_mult_53(244);
partial_product_2(245) <= temp_mult_53(245);
partial_product_2(246) <= temp_mult_53(246);
partial_product_2(247) <= temp_mult_53(247);
partial_product_2(248) <= temp_mult_53(248);
partial_product_2(249) <= temp_mult_53(249);
partial_product_2(250) <= temp_mult_53(250);
partial_product_2(251) <= temp_mult_53(251);
partial_product_2(252) <= temp_mult_53(252);
partial_product_2(253) <= temp_mult_53(253);
partial_product_2(254) <= temp_mult_53(254);
partial_product_2(255) <= temp_mult_53(255);
partial_product_2(256) <= temp_mult_53(256);
partial_product_2(257) <= temp_mult_53(257);
partial_product_2(258) <= temp_mult_53(258);
partial_product_2(259) <= temp_mult_53(259);
partial_product_2(260) <= temp_mult_53(260);
partial_product_2(261) <= temp_mult_53(261);
partial_product_2(262) <= temp_mult_53(262);
partial_product_2(263) <= temp_mult_53(263);
partial_product_2(264) <= temp_mult_53(264);
partial_product_2(265) <= temp_mult_53(265);
partial_product_2(266) <= temp_mult_53(266);
partial_product_2(267) <= temp_mult_53(267);
partial_product_2(268) <= temp_mult_53(268);
partial_product_2(269) <= temp_mult_53(269);
partial_product_2(270) <= temp_mult_62(270);
partial_product_2(271) <= temp_mult_62(271);
partial_product_2(272) <= temp_mult_62(272);
partial_product_2(273) <= temp_mult_62(273);
partial_product_2(274) <= temp_mult_62(274);
partial_product_2(275) <= temp_mult_62(275);
partial_product_2(276) <= temp_mult_62(276);
partial_product_2(277) <= temp_mult_62(277);
partial_product_2(278) <= temp_mult_62(278);
partial_product_2(279) <= temp_mult_62(279);
partial_product_2(280) <= temp_mult_62(280);
partial_product_2(281) <= temp_mult_62(281);
partial_product_2(282) <= temp_mult_62(282);
partial_product_2(283) <= temp_mult_62(283);
partial_product_2(284) <= temp_mult_62(284);
partial_product_2(285) <= temp_mult_62(285);
partial_product_2(286) <= temp_mult_62(286);
partial_product_2(287) <= temp_mult_62(287);
partial_product_2(288) <= temp_mult_62(288);
partial_product_2(289) <= temp_mult_62(289);
partial_product_2(290) <= temp_mult_62(290);
partial_product_2(291) <= temp_mult_62(291);
partial_product_2(292) <= temp_mult_62(292);
partial_product_2(293) <= temp_mult_62(293);
partial_product_2(294) <= temp_mult_62(294);
partial_product_2(295) <= temp_mult_62(295);
partial_product_2(296) <= temp_mult_62(296);
partial_product_2(297) <= temp_mult_62(297);
partial_product_2(298) <= temp_mult_62(298);
partial_product_2(299) <= temp_mult_62(299);
partial_product_2(300) <= temp_mult_62(300);
partial_product_2(301) <= temp_mult_62(301);
partial_product_2(302) <= temp_mult_62(302);
partial_product_2(303) <= temp_mult_62(303);
partial_product_2(304) <= temp_mult_62(304);
partial_product_2(305) <= temp_mult_62(305);
partial_product_2(306) <= temp_mult_62(306);
partial_product_2(307) <= temp_mult_62(307);
partial_product_2(308) <= temp_mult_62(308);
partial_product_2(309) <= temp_mult_62(309);
partial_product_2(310) <= temp_mult_62(310);
partial_product_2(311) <= temp_mult_71(311);
partial_product_2(312) <= temp_mult_71(312);
partial_product_2(313) <= temp_mult_71(313);
partial_product_2(314) <= temp_mult_71(314);
partial_product_2(315) <= temp_mult_71(315);
partial_product_2(316) <= temp_mult_71(316);
partial_product_2(317) <= temp_mult_71(317);
partial_product_2(318) <= temp_mult_71(318);
partial_product_2(319) <= temp_mult_71(319);
partial_product_2(320) <= temp_mult_71(320);
partial_product_2(321) <= temp_mult_71(321);
partial_product_2(322) <= temp_mult_71(322);
partial_product_2(323) <= temp_mult_71(323);
partial_product_2(324) <= temp_mult_71(324);
partial_product_2(325) <= temp_mult_71(325);
partial_product_2(326) <= temp_mult_71(326);
partial_product_2(327) <= temp_mult_71(327);
partial_product_2(328) <= temp_mult_71(328);
partial_product_2(329) <= temp_mult_71(329);
partial_product_2(330) <= temp_mult_71(330);
partial_product_2(331) <= temp_mult_71(331);
partial_product_2(332) <= temp_mult_71(332);
partial_product_2(333) <= temp_mult_71(333);
partial_product_2(334) <= temp_mult_71(334);
partial_product_2(335) <= temp_mult_71(335);
partial_product_2(336) <= temp_mult_71(336);
partial_product_2(337) <= temp_mult_71(337);
partial_product_2(338) <= temp_mult_71(338);
partial_product_2(339) <= temp_mult_71(339);
partial_product_2(340) <= temp_mult_71(340);
partial_product_2(341) <= temp_mult_71(341);
partial_product_2(342) <= temp_mult_71(342);
partial_product_2(343) <= temp_mult_71(343);
partial_product_2(344) <= temp_mult_71(344);
partial_product_2(345) <= temp_mult_71(345);
partial_product_2(346) <= temp_mult_71(346);
partial_product_2(347) <= temp_mult_71(347);
partial_product_2(348) <= temp_mult_71(348);
partial_product_2(349) <= temp_mult_71(349);
partial_product_2(350) <= temp_mult_71(350);
partial_product_2(351) <= temp_mult_71(351);
partial_product_2(352) <= temp_mult_124(352);
partial_product_2(353) <= temp_mult_124(353);
partial_product_2(354) <= temp_mult_124(354);
partial_product_2(355) <= temp_mult_124(355);
partial_product_2(356) <= temp_mult_124(356);
partial_product_2(357) <= temp_mult_124(357);
partial_product_2(358) <= temp_mult_124(358);
partial_product_2(359) <= temp_mult_124(359);
partial_product_2(360) <= temp_mult_124(360);
partial_product_2(361) <= temp_mult_124(361);
partial_product_2(362) <= temp_mult_124(362);
partial_product_2(363) <= temp_mult_124(363);
partial_product_2(364) <= temp_mult_124(364);
partial_product_2(365) <= temp_mult_124(365);
partial_product_2(366) <= temp_mult_124(366);
partial_product_2(367) <= temp_mult_124(367);
partial_product_2(368) <= temp_mult_124(368);
partial_product_2(369) <= temp_mult_124(369);
partial_product_2(370) <= temp_mult_124(370);
partial_product_2(371) <= temp_mult_124(371);
partial_product_2(372) <= temp_mult_124(372);
partial_product_2(373) <= temp_mult_124(373);
partial_product_2(374) <= temp_mult_124(374);
partial_product_2(375) <= temp_mult_124(375);
partial_product_2(376) <= temp_mult_124(376);
partial_product_2(377) <= temp_mult_124(377);
partial_product_2(378) <= temp_mult_124(378);
partial_product_2(379) <= temp_mult_124(379);
partial_product_2(380) <= temp_mult_124(380);
partial_product_2(381) <= temp_mult_124(381);
partial_product_2(382) <= temp_mult_124(382);
partial_product_2(383) <= temp_mult_124(383);
partial_product_2(384) <= temp_mult_124(384);
partial_product_2(385) <= temp_mult_124(385);
partial_product_2(386) <= temp_mult_124(386);
partial_product_2(387) <= temp_mult_124(387);
partial_product_2(388) <= temp_mult_124(388);
partial_product_2(389) <= temp_mult_124(389);
partial_product_2(390) <= temp_mult_124(390);
partial_product_2(391) <= temp_mult_124(391);
partial_product_2(392) <= temp_mult_124(392);
partial_product_2(393) <= '0';
partial_product_2(394) <= '0';
partial_product_2(395) <= '0';
partial_product_2(396) <= temp_mult_143(396);
partial_product_2(397) <= temp_mult_143(397);
partial_product_2(398) <= temp_mult_143(398);
partial_product_2(399) <= temp_mult_143(399);
partial_product_2(400) <= temp_mult_143(400);
partial_product_2(401) <= temp_mult_143(401);
partial_product_2(402) <= temp_mult_143(402);
partial_product_2(403) <= temp_mult_143(403);
partial_product_2(404) <= temp_mult_143(404);
partial_product_2(405) <= temp_mult_143(405);
partial_product_2(406) <= temp_mult_143(406);
partial_product_2(407) <= temp_mult_143(407);
partial_product_2(408) <= temp_mult_143(408);
partial_product_2(409) <= temp_mult_143(409);
partial_product_2(410) <= temp_mult_143(410);
partial_product_2(411) <= temp_mult_143(411);
partial_product_2(412) <= temp_mult_143(412);
partial_product_2(413) <= temp_mult_143(413);
partial_product_2(414) <= temp_mult_143(414);
partial_product_2(415) <= temp_mult_143(415);
partial_product_2(416) <= temp_mult_143(416);
partial_product_2(417) <= temp_mult_143(417);
partial_product_2(418) <= temp_mult_143(418);
partial_product_2(419) <= temp_mult_143(419);
partial_product_2(420) <= temp_mult_143(420);
partial_product_2(421) <= temp_mult_143(421);
partial_product_2(422) <= temp_mult_143(422);
partial_product_2(423) <= temp_mult_143(423);
partial_product_2(424) <= temp_mult_143(424);
partial_product_2(425) <= temp_mult_143(425);
partial_product_2(426) <= temp_mult_143(426);
partial_product_2(427) <= temp_mult_143(427);
partial_product_2(428) <= temp_mult_143(428);
partial_product_2(429) <= temp_mult_143(429);
partial_product_2(430) <= temp_mult_143(430);
partial_product_2(431) <= temp_mult_143(431);
partial_product_2(432) <= temp_mult_143(432);
partial_product_2(433) <= temp_mult_143(433);
partial_product_2(434) <= temp_mult_143(434);
partial_product_2(435) <= temp_mult_143(435);
partial_product_2(436) <= temp_mult_143(436);
partial_product_2(437) <= temp_mult_149(437);
partial_product_2(438) <= temp_mult_149(438);
partial_product_2(439) <= temp_mult_149(439);
partial_product_2(440) <= temp_mult_149(440);
partial_product_2(441) <= temp_mult_149(441);
partial_product_2(442) <= temp_mult_149(442);
partial_product_2(443) <= temp_mult_149(443);
partial_product_2(444) <= temp_mult_149(444);
partial_product_2(445) <= temp_mult_149(445);
partial_product_2(446) <= temp_mult_149(446);
partial_product_2(447) <= temp_mult_149(447);
partial_product_2(448) <= temp_mult_149(448);
partial_product_2(449) <= temp_mult_149(449);
partial_product_2(450) <= temp_mult_149(450);
partial_product_2(451) <= temp_mult_149(451);
partial_product_2(452) <= temp_mult_149(452);
partial_product_2(453) <= temp_mult_149(453);
partial_product_2(454) <= temp_mult_149(454);
partial_product_2(455) <= temp_mult_149(455);
partial_product_2(456) <= temp_mult_149(456);
partial_product_2(457) <= temp_mult_149(457);
partial_product_2(458) <= temp_mult_149(458);
partial_product_2(459) <= temp_mult_149(459);
partial_product_2(460) <= temp_mult_149(460);
partial_product_2(461) <= temp_mult_149(461);
partial_product_2(462) <= temp_mult_149(462);
partial_product_2(463) <= temp_mult_149(463);
partial_product_2(464) <= temp_mult_149(464);
partial_product_2(465) <= temp_mult_149(465);
partial_product_2(466) <= temp_mult_149(466);
partial_product_2(467) <= temp_mult_149(467);
partial_product_2(468) <= temp_mult_149(468);
partial_product_2(469) <= temp_mult_149(469);
partial_product_2(470) <= temp_mult_149(470);
partial_product_2(471) <= temp_mult_149(471);
partial_product_2(472) <= temp_mult_149(472);
partial_product_2(473) <= temp_mult_149(473);
partial_product_2(474) <= temp_mult_149(474);
partial_product_2(475) <= temp_mult_149(475);
partial_product_2(476) <= temp_mult_149(476);
partial_product_2(477) <= temp_mult_149(477);
partial_product_2(478) <= '0';
partial_product_2(479) <= '0';
partial_product_2(480) <= '0';
partial_product_2(481) <= '0';
partial_product_2(482) <= '0';
partial_product_2(483) <= '0';
partial_product_2(484) <= '0';
partial_product_2(485) <= '0';
partial_product_2(486) <= '0';
partial_product_2(487) <= '0';
partial_product_2(488) <= '0';
partial_product_2(489) <= '0';
partial_product_2(490) <= '0';
partial_product_2(491) <= '0';
partial_product_2(492) <= '0';
partial_product_2(493) <= '0';
partial_product_2(494) <= '0';
partial_product_2(495) <= '0';
partial_product_2(496) <= '0';
partial_product_2(497) <= '0';
partial_product_2(498) <= '0';
partial_product_2(499) <= '0';
partial_product_2(500) <= '0';
partial_product_2(501) <= '0';
partial_product_2(502) <= '0';
partial_product_2(503) <= '0';
partial_product_2(504) <= '0';
partial_product_2(505) <= '0';
partial_product_2(506) <= '0';
partial_product_2(507) <= '0';
partial_product_2(508) <= '0';
partial_product_2(509) <= '0';
partial_product_2(510) <= '0';
partial_product_2(511) <= '0';
partial_product_2(512) <= '0';
partial_product_3(0) <= '0';
partial_product_3(1) <= '0';
partial_product_3(2) <= '0';
partial_product_3(3) <= '0';
partial_product_3(4) <= '0';
partial_product_3(5) <= '0';
partial_product_3(6) <= '0';
partial_product_3(7) <= '0';
partial_product_3(8) <= '0';
partial_product_3(9) <= '0';
partial_product_3(10) <= '0';
partial_product_3(11) <= '0';
partial_product_3(12) <= '0';
partial_product_3(13) <= '0';
partial_product_3(14) <= '0';
partial_product_3(15) <= '0';
partial_product_3(16) <= '0';
partial_product_3(17) <= '0';
partial_product_3(18) <= '0';
partial_product_3(19) <= '0';
partial_product_3(20) <= '0';
partial_product_3(21) <= '0';
partial_product_3(22) <= '0';
partial_product_3(23) <= '0';
partial_product_3(24) <= '0';
partial_product_3(25) <= '0';
partial_product_3(26) <= '0';
partial_product_3(27) <= '0';
partial_product_3(28) <= '0';
partial_product_3(29) <= '0';
partial_product_3(30) <= '0';
partial_product_3(31) <= '0';
partial_product_3(32) <= '0';
partial_product_3(33) <= '0';
partial_product_3(34) <= temp_mult_10(34);
partial_product_3(35) <= temp_mult_10(35);
partial_product_3(36) <= temp_mult_10(36);
partial_product_3(37) <= temp_mult_10(37);
partial_product_3(38) <= temp_mult_10(38);
partial_product_3(39) <= temp_mult_10(39);
partial_product_3(40) <= temp_mult_10(40);
partial_product_3(41) <= temp_mult_10(41);
partial_product_3(42) <= temp_mult_10(42);
partial_product_3(43) <= temp_mult_10(43);
partial_product_3(44) <= temp_mult_10(44);
partial_product_3(45) <= temp_mult_10(45);
partial_product_3(46) <= temp_mult_10(46);
partial_product_3(47) <= temp_mult_10(47);
partial_product_3(48) <= temp_mult_10(48);
partial_product_3(49) <= temp_mult_10(49);
partial_product_3(50) <= temp_mult_10(50);
partial_product_3(51) <= temp_mult_10(51);
partial_product_3(52) <= temp_mult_10(52);
partial_product_3(53) <= temp_mult_10(53);
partial_product_3(54) <= temp_mult_10(54);
partial_product_3(55) <= temp_mult_10(55);
partial_product_3(56) <= temp_mult_10(56);
partial_product_3(57) <= temp_mult_10(57);
partial_product_3(58) <= temp_mult_10(58);
partial_product_3(59) <= temp_mult_10(59);
partial_product_3(60) <= temp_mult_10(60);
partial_product_3(61) <= temp_mult_10(61);
partial_product_3(62) <= temp_mult_10(62);
partial_product_3(63) <= temp_mult_10(63);
partial_product_3(64) <= temp_mult_10(64);
partial_product_3(65) <= temp_mult_10(65);
partial_product_3(66) <= temp_mult_10(66);
partial_product_3(67) <= temp_mult_10(67);
partial_product_3(68) <= temp_mult_10(68);
partial_product_3(69) <= temp_mult_10(69);
partial_product_3(70) <= temp_mult_10(70);
partial_product_3(71) <= temp_mult_10(71);
partial_product_3(72) <= temp_mult_10(72);
partial_product_3(73) <= temp_mult_10(73);
partial_product_3(74) <= temp_mult_10(74);
partial_product_3(75) <= temp_mult_16(75);
partial_product_3(76) <= temp_mult_16(76);
partial_product_3(77) <= temp_mult_16(77);
partial_product_3(78) <= temp_mult_16(78);
partial_product_3(79) <= temp_mult_16(79);
partial_product_3(80) <= temp_mult_16(80);
partial_product_3(81) <= temp_mult_16(81);
partial_product_3(82) <= temp_mult_16(82);
partial_product_3(83) <= temp_mult_16(83);
partial_product_3(84) <= temp_mult_16(84);
partial_product_3(85) <= temp_mult_16(85);
partial_product_3(86) <= temp_mult_16(86);
partial_product_3(87) <= temp_mult_16(87);
partial_product_3(88) <= temp_mult_16(88);
partial_product_3(89) <= temp_mult_16(89);
partial_product_3(90) <= temp_mult_16(90);
partial_product_3(91) <= temp_mult_16(91);
partial_product_3(92) <= temp_mult_16(92);
partial_product_3(93) <= temp_mult_16(93);
partial_product_3(94) <= temp_mult_16(94);
partial_product_3(95) <= temp_mult_16(95);
partial_product_3(96) <= temp_mult_16(96);
partial_product_3(97) <= temp_mult_16(97);
partial_product_3(98) <= temp_mult_16(98);
partial_product_3(99) <= temp_mult_16(99);
partial_product_3(100) <= temp_mult_16(100);
partial_product_3(101) <= temp_mult_16(101);
partial_product_3(102) <= temp_mult_16(102);
partial_product_3(103) <= temp_mult_16(103);
partial_product_3(104) <= temp_mult_16(104);
partial_product_3(105) <= temp_mult_16(105);
partial_product_3(106) <= temp_mult_16(106);
partial_product_3(107) <= temp_mult_16(107);
partial_product_3(108) <= temp_mult_16(108);
partial_product_3(109) <= temp_mult_16(109);
partial_product_3(110) <= temp_mult_16(110);
partial_product_3(111) <= temp_mult_16(111);
partial_product_3(112) <= temp_mult_16(112);
partial_product_3(113) <= temp_mult_16(113);
partial_product_3(114) <= temp_mult_16(114);
partial_product_3(115) <= temp_mult_16(115);
partial_product_3(116) <= temp_mult_22(116);
partial_product_3(117) <= temp_mult_22(117);
partial_product_3(118) <= temp_mult_22(118);
partial_product_3(119) <= temp_mult_22(119);
partial_product_3(120) <= temp_mult_22(120);
partial_product_3(121) <= temp_mult_22(121);
partial_product_3(122) <= temp_mult_22(122);
partial_product_3(123) <= temp_mult_22(123);
partial_product_3(124) <= temp_mult_22(124);
partial_product_3(125) <= temp_mult_22(125);
partial_product_3(126) <= temp_mult_22(126);
partial_product_3(127) <= temp_mult_22(127);
partial_product_3(128) <= temp_mult_22(128);
partial_product_3(129) <= temp_mult_22(129);
partial_product_3(130) <= temp_mult_22(130);
partial_product_3(131) <= temp_mult_22(131);
partial_product_3(132) <= temp_mult_22(132);
partial_product_3(133) <= temp_mult_22(133);
partial_product_3(134) <= temp_mult_22(134);
partial_product_3(135) <= temp_mult_22(135);
partial_product_3(136) <= temp_mult_22(136);
partial_product_3(137) <= temp_mult_22(137);
partial_product_3(138) <= temp_mult_22(138);
partial_product_3(139) <= temp_mult_22(139);
partial_product_3(140) <= temp_mult_22(140);
partial_product_3(141) <= temp_mult_22(141);
partial_product_3(142) <= temp_mult_22(142);
partial_product_3(143) <= temp_mult_22(143);
partial_product_3(144) <= temp_mult_22(144);
partial_product_3(145) <= temp_mult_22(145);
partial_product_3(146) <= temp_mult_22(146);
partial_product_3(147) <= temp_mult_22(147);
partial_product_3(148) <= temp_mult_22(148);
partial_product_3(149) <= temp_mult_22(149);
partial_product_3(150) <= temp_mult_22(150);
partial_product_3(151) <= temp_mult_22(151);
partial_product_3(152) <= temp_mult_22(152);
partial_product_3(153) <= temp_mult_22(153);
partial_product_3(154) <= temp_mult_22(154);
partial_product_3(155) <= temp_mult_22(155);
partial_product_3(156) <= temp_mult_22(156);
partial_product_3(157) <= temp_mult_28(157);
partial_product_3(158) <= temp_mult_28(158);
partial_product_3(159) <= temp_mult_28(159);
partial_product_3(160) <= temp_mult_28(160);
partial_product_3(161) <= temp_mult_28(161);
partial_product_3(162) <= temp_mult_28(162);
partial_product_3(163) <= temp_mult_28(163);
partial_product_3(164) <= temp_mult_28(164);
partial_product_3(165) <= temp_mult_28(165);
partial_product_3(166) <= temp_mult_28(166);
partial_product_3(167) <= temp_mult_28(167);
partial_product_3(168) <= temp_mult_28(168);
partial_product_3(169) <= temp_mult_28(169);
partial_product_3(170) <= temp_mult_28(170);
partial_product_3(171) <= temp_mult_28(171);
partial_product_3(172) <= temp_mult_28(172);
partial_product_3(173) <= temp_mult_28(173);
partial_product_3(174) <= temp_mult_28(174);
partial_product_3(175) <= temp_mult_28(175);
partial_product_3(176) <= temp_mult_28(176);
partial_product_3(177) <= temp_mult_28(177);
partial_product_3(178) <= temp_mult_28(178);
partial_product_3(179) <= temp_mult_28(179);
partial_product_3(180) <= temp_mult_28(180);
partial_product_3(181) <= temp_mult_28(181);
partial_product_3(182) <= temp_mult_28(182);
partial_product_3(183) <= temp_mult_28(183);
partial_product_3(184) <= temp_mult_28(184);
partial_product_3(185) <= temp_mult_28(185);
partial_product_3(186) <= temp_mult_28(186);
partial_product_3(187) <= temp_mult_28(187);
partial_product_3(188) <= temp_mult_28(188);
partial_product_3(189) <= temp_mult_28(189);
partial_product_3(190) <= temp_mult_28(190);
partial_product_3(191) <= temp_mult_28(191);
partial_product_3(192) <= temp_mult_28(192);
partial_product_3(193) <= temp_mult_28(193);
partial_product_3(194) <= temp_mult_28(194);
partial_product_3(195) <= temp_mult_28(195);
partial_product_3(196) <= temp_mult_28(196);
partial_product_3(197) <= temp_mult_28(197);
partial_product_3(198) <= temp_mult_34(198);
partial_product_3(199) <= temp_mult_34(199);
partial_product_3(200) <= temp_mult_34(200);
partial_product_3(201) <= temp_mult_34(201);
partial_product_3(202) <= temp_mult_34(202);
partial_product_3(203) <= temp_mult_34(203);
partial_product_3(204) <= temp_mult_34(204);
partial_product_3(205) <= temp_mult_34(205);
partial_product_3(206) <= temp_mult_34(206);
partial_product_3(207) <= temp_mult_34(207);
partial_product_3(208) <= temp_mult_34(208);
partial_product_3(209) <= temp_mult_34(209);
partial_product_3(210) <= temp_mult_34(210);
partial_product_3(211) <= temp_mult_34(211);
partial_product_3(212) <= temp_mult_34(212);
partial_product_3(213) <= temp_mult_34(213);
partial_product_3(214) <= temp_mult_34(214);
partial_product_3(215) <= temp_mult_34(215);
partial_product_3(216) <= temp_mult_34(216);
partial_product_3(217) <= temp_mult_34(217);
partial_product_3(218) <= temp_mult_34(218);
partial_product_3(219) <= temp_mult_34(219);
partial_product_3(220) <= temp_mult_34(220);
partial_product_3(221) <= temp_mult_34(221);
partial_product_3(222) <= temp_mult_34(222);
partial_product_3(223) <= temp_mult_34(223);
partial_product_3(224) <= temp_mult_34(224);
partial_product_3(225) <= temp_mult_34(225);
partial_product_3(226) <= temp_mult_34(226);
partial_product_3(227) <= temp_mult_34(227);
partial_product_3(228) <= temp_mult_34(228);
partial_product_3(229) <= temp_mult_34(229);
partial_product_3(230) <= temp_mult_34(230);
partial_product_3(231) <= temp_mult_34(231);
partial_product_3(232) <= temp_mult_34(232);
partial_product_3(233) <= temp_mult_34(233);
partial_product_3(234) <= temp_mult_34(234);
partial_product_3(235) <= temp_mult_34(235);
partial_product_3(236) <= temp_mult_34(236);
partial_product_3(237) <= temp_mult_34(237);
partial_product_3(238) <= temp_mult_34(238);
partial_product_3(239) <= temp_mult_47(239);
partial_product_3(240) <= temp_mult_47(240);
partial_product_3(241) <= temp_mult_47(241);
partial_product_3(242) <= temp_mult_47(242);
partial_product_3(243) <= temp_mult_47(243);
partial_product_3(244) <= temp_mult_47(244);
partial_product_3(245) <= temp_mult_47(245);
partial_product_3(246) <= temp_mult_47(246);
partial_product_3(247) <= temp_mult_47(247);
partial_product_3(248) <= temp_mult_47(248);
partial_product_3(249) <= temp_mult_47(249);
partial_product_3(250) <= temp_mult_47(250);
partial_product_3(251) <= temp_mult_47(251);
partial_product_3(252) <= temp_mult_47(252);
partial_product_3(253) <= temp_mult_47(253);
partial_product_3(254) <= temp_mult_47(254);
partial_product_3(255) <= temp_mult_47(255);
partial_product_3(256) <= temp_mult_47(256);
partial_product_3(257) <= temp_mult_47(257);
partial_product_3(258) <= temp_mult_47(258);
partial_product_3(259) <= temp_mult_47(259);
partial_product_3(260) <= temp_mult_47(260);
partial_product_3(261) <= temp_mult_47(261);
partial_product_3(262) <= temp_mult_47(262);
partial_product_3(263) <= temp_mult_47(263);
partial_product_3(264) <= temp_mult_47(264);
partial_product_3(265) <= temp_mult_47(265);
partial_product_3(266) <= temp_mult_47(266);
partial_product_3(267) <= temp_mult_47(267);
partial_product_3(268) <= temp_mult_47(268);
partial_product_3(269) <= temp_mult_47(269);
partial_product_3(270) <= temp_mult_47(270);
partial_product_3(271) <= temp_mult_47(271);
partial_product_3(272) <= temp_mult_47(272);
partial_product_3(273) <= temp_mult_47(273);
partial_product_3(274) <= temp_mult_47(274);
partial_product_3(275) <= temp_mult_47(275);
partial_product_3(276) <= temp_mult_47(276);
partial_product_3(277) <= temp_mult_47(277);
partial_product_3(278) <= temp_mult_47(278);
partial_product_3(279) <= temp_mult_47(279);
partial_product_3(280) <= temp_mult_121(280);
partial_product_3(281) <= temp_mult_121(281);
partial_product_3(282) <= temp_mult_121(282);
partial_product_3(283) <= temp_mult_121(283);
partial_product_3(284) <= temp_mult_121(284);
partial_product_3(285) <= temp_mult_121(285);
partial_product_3(286) <= temp_mult_121(286);
partial_product_3(287) <= temp_mult_121(287);
partial_product_3(288) <= temp_mult_121(288);
partial_product_3(289) <= temp_mult_121(289);
partial_product_3(290) <= temp_mult_121(290);
partial_product_3(291) <= temp_mult_121(291);
partial_product_3(292) <= temp_mult_121(292);
partial_product_3(293) <= temp_mult_121(293);
partial_product_3(294) <= temp_mult_121(294);
partial_product_3(295) <= temp_mult_121(295);
partial_product_3(296) <= temp_mult_121(296);
partial_product_3(297) <= temp_mult_121(297);
partial_product_3(298) <= temp_mult_121(298);
partial_product_3(299) <= temp_mult_121(299);
partial_product_3(300) <= temp_mult_121(300);
partial_product_3(301) <= temp_mult_121(301);
partial_product_3(302) <= temp_mult_121(302);
partial_product_3(303) <= temp_mult_121(303);
partial_product_3(304) <= temp_mult_121(304);
partial_product_3(305) <= temp_mult_121(305);
partial_product_3(306) <= temp_mult_121(306);
partial_product_3(307) <= temp_mult_121(307);
partial_product_3(308) <= temp_mult_121(308);
partial_product_3(309) <= temp_mult_121(309);
partial_product_3(310) <= temp_mult_121(310);
partial_product_3(311) <= temp_mult_121(311);
partial_product_3(312) <= temp_mult_121(312);
partial_product_3(313) <= temp_mult_121(313);
partial_product_3(314) <= temp_mult_121(314);
partial_product_3(315) <= temp_mult_121(315);
partial_product_3(316) <= temp_mult_121(316);
partial_product_3(317) <= temp_mult_121(317);
partial_product_3(318) <= temp_mult_121(318);
partial_product_3(319) <= temp_mult_121(319);
partial_product_3(320) <= temp_mult_121(320);
partial_product_3(321) <= temp_mult_127(321);
partial_product_3(322) <= temp_mult_127(322);
partial_product_3(323) <= temp_mult_127(323);
partial_product_3(324) <= temp_mult_127(324);
partial_product_3(325) <= temp_mult_127(325);
partial_product_3(326) <= temp_mult_127(326);
partial_product_3(327) <= temp_mult_127(327);
partial_product_3(328) <= temp_mult_127(328);
partial_product_3(329) <= temp_mult_127(329);
partial_product_3(330) <= temp_mult_127(330);
partial_product_3(331) <= temp_mult_127(331);
partial_product_3(332) <= temp_mult_127(332);
partial_product_3(333) <= temp_mult_127(333);
partial_product_3(334) <= temp_mult_127(334);
partial_product_3(335) <= temp_mult_127(335);
partial_product_3(336) <= temp_mult_127(336);
partial_product_3(337) <= temp_mult_127(337);
partial_product_3(338) <= temp_mult_127(338);
partial_product_3(339) <= temp_mult_127(339);
partial_product_3(340) <= temp_mult_127(340);
partial_product_3(341) <= temp_mult_127(341);
partial_product_3(342) <= temp_mult_127(342);
partial_product_3(343) <= temp_mult_127(343);
partial_product_3(344) <= temp_mult_127(344);
partial_product_3(345) <= temp_mult_127(345);
partial_product_3(346) <= temp_mult_127(346);
partial_product_3(347) <= temp_mult_127(347);
partial_product_3(348) <= temp_mult_127(348);
partial_product_3(349) <= temp_mult_127(349);
partial_product_3(350) <= temp_mult_127(350);
partial_product_3(351) <= temp_mult_127(351);
partial_product_3(352) <= temp_mult_127(352);
partial_product_3(353) <= temp_mult_127(353);
partial_product_3(354) <= temp_mult_127(354);
partial_product_3(355) <= temp_mult_127(355);
partial_product_3(356) <= temp_mult_127(356);
partial_product_3(357) <= temp_mult_127(357);
partial_product_3(358) <= temp_mult_127(358);
partial_product_3(359) <= temp_mult_127(359);
partial_product_3(360) <= temp_mult_127(360);
partial_product_3(361) <= temp_mult_127(361);
partial_product_3(362) <= temp_mult_133(362);
partial_product_3(363) <= temp_mult_133(363);
partial_product_3(364) <= temp_mult_133(364);
partial_product_3(365) <= temp_mult_133(365);
partial_product_3(366) <= temp_mult_133(366);
partial_product_3(367) <= temp_mult_133(367);
partial_product_3(368) <= temp_mult_133(368);
partial_product_3(369) <= temp_mult_133(369);
partial_product_3(370) <= temp_mult_133(370);
partial_product_3(371) <= temp_mult_133(371);
partial_product_3(372) <= temp_mult_133(372);
partial_product_3(373) <= temp_mult_133(373);
partial_product_3(374) <= temp_mult_133(374);
partial_product_3(375) <= temp_mult_133(375);
partial_product_3(376) <= temp_mult_133(376);
partial_product_3(377) <= temp_mult_133(377);
partial_product_3(378) <= temp_mult_133(378);
partial_product_3(379) <= temp_mult_133(379);
partial_product_3(380) <= temp_mult_133(380);
partial_product_3(381) <= temp_mult_133(381);
partial_product_3(382) <= temp_mult_133(382);
partial_product_3(383) <= temp_mult_133(383);
partial_product_3(384) <= temp_mult_133(384);
partial_product_3(385) <= temp_mult_133(385);
partial_product_3(386) <= temp_mult_133(386);
partial_product_3(387) <= temp_mult_133(387);
partial_product_3(388) <= temp_mult_133(388);
partial_product_3(389) <= temp_mult_133(389);
partial_product_3(390) <= temp_mult_133(390);
partial_product_3(391) <= temp_mult_133(391);
partial_product_3(392) <= temp_mult_133(392);
partial_product_3(393) <= temp_mult_133(393);
partial_product_3(394) <= temp_mult_133(394);
partial_product_3(395) <= temp_mult_133(395);
partial_product_3(396) <= temp_mult_133(396);
partial_product_3(397) <= temp_mult_133(397);
partial_product_3(398) <= temp_mult_133(398);
partial_product_3(399) <= temp_mult_133(399);
partial_product_3(400) <= temp_mult_133(400);
partial_product_3(401) <= temp_mult_133(401);
partial_product_3(402) <= temp_mult_133(402);
partial_product_3(403) <= temp_mult_139(403);
partial_product_3(404) <= temp_mult_139(404);
partial_product_3(405) <= temp_mult_139(405);
partial_product_3(406) <= temp_mult_139(406);
partial_product_3(407) <= temp_mult_139(407);
partial_product_3(408) <= temp_mult_139(408);
partial_product_3(409) <= temp_mult_139(409);
partial_product_3(410) <= temp_mult_139(410);
partial_product_3(411) <= temp_mult_139(411);
partial_product_3(412) <= temp_mult_139(412);
partial_product_3(413) <= temp_mult_139(413);
partial_product_3(414) <= temp_mult_139(414);
partial_product_3(415) <= temp_mult_139(415);
partial_product_3(416) <= temp_mult_139(416);
partial_product_3(417) <= temp_mult_139(417);
partial_product_3(418) <= temp_mult_139(418);
partial_product_3(419) <= temp_mult_139(419);
partial_product_3(420) <= temp_mult_139(420);
partial_product_3(421) <= temp_mult_139(421);
partial_product_3(422) <= temp_mult_139(422);
partial_product_3(423) <= temp_mult_139(423);
partial_product_3(424) <= temp_mult_139(424);
partial_product_3(425) <= temp_mult_139(425);
partial_product_3(426) <= temp_mult_139(426);
partial_product_3(427) <= temp_mult_139(427);
partial_product_3(428) <= temp_mult_139(428);
partial_product_3(429) <= temp_mult_139(429);
partial_product_3(430) <= temp_mult_139(430);
partial_product_3(431) <= temp_mult_139(431);
partial_product_3(432) <= temp_mult_139(432);
partial_product_3(433) <= temp_mult_139(433);
partial_product_3(434) <= temp_mult_139(434);
partial_product_3(435) <= temp_mult_139(435);
partial_product_3(436) <= temp_mult_139(436);
partial_product_3(437) <= temp_mult_139(437);
partial_product_3(438) <= temp_mult_139(438);
partial_product_3(439) <= temp_mult_139(439);
partial_product_3(440) <= temp_mult_139(440);
partial_product_3(441) <= temp_mult_139(441);
partial_product_3(442) <= temp_mult_139(442);
partial_product_3(443) <= temp_mult_139(443);
partial_product_3(444) <= '0';
partial_product_3(445) <= '0';
partial_product_3(446) <= '0';
partial_product_3(447) <= temp_mult_158(447);
partial_product_3(448) <= temp_mult_158(448);
partial_product_3(449) <= temp_mult_158(449);
partial_product_3(450) <= temp_mult_158(450);
partial_product_3(451) <= temp_mult_158(451);
partial_product_3(452) <= temp_mult_158(452);
partial_product_3(453) <= temp_mult_158(453);
partial_product_3(454) <= temp_mult_158(454);
partial_product_3(455) <= temp_mult_158(455);
partial_product_3(456) <= temp_mult_158(456);
partial_product_3(457) <= temp_mult_158(457);
partial_product_3(458) <= temp_mult_158(458);
partial_product_3(459) <= temp_mult_158(459);
partial_product_3(460) <= temp_mult_158(460);
partial_product_3(461) <= temp_mult_158(461);
partial_product_3(462) <= temp_mult_158(462);
partial_product_3(463) <= temp_mult_158(463);
partial_product_3(464) <= temp_mult_158(464);
partial_product_3(465) <= temp_mult_158(465);
partial_product_3(466) <= temp_mult_158(466);
partial_product_3(467) <= temp_mult_158(467);
partial_product_3(468) <= temp_mult_158(468);
partial_product_3(469) <= temp_mult_158(469);
partial_product_3(470) <= temp_mult_158(470);
partial_product_3(471) <= temp_mult_158(471);
partial_product_3(472) <= temp_mult_158(472);
partial_product_3(473) <= temp_mult_158(473);
partial_product_3(474) <= temp_mult_158(474);
partial_product_3(475) <= temp_mult_158(475);
partial_product_3(476) <= temp_mult_158(476);
partial_product_3(477) <= temp_mult_158(477);
partial_product_3(478) <= temp_mult_158(478);
partial_product_3(479) <= temp_mult_158(479);
partial_product_3(480) <= temp_mult_158(480);
partial_product_3(481) <= temp_mult_158(481);
partial_product_3(482) <= temp_mult_158(482);
partial_product_3(483) <= temp_mult_158(483);
partial_product_3(484) <= temp_mult_158(484);
partial_product_3(485) <= temp_mult_158(485);
partial_product_3(486) <= temp_mult_158(486);
partial_product_3(487) <= temp_mult_158(487);
partial_product_3(488) <= '0';
partial_product_3(489) <= '0';
partial_product_3(490) <= '0';
partial_product_3(491) <= '0';
partial_product_3(492) <= '0';
partial_product_3(493) <= '0';
partial_product_3(494) <= '0';
partial_product_3(495) <= '0';
partial_product_3(496) <= '0';
partial_product_3(497) <= '0';
partial_product_3(498) <= '0';
partial_product_3(499) <= '0';
partial_product_3(500) <= '0';
partial_product_3(501) <= '0';
partial_product_3(502) <= '0';
partial_product_3(503) <= '0';
partial_product_3(504) <= '0';
partial_product_3(505) <= '0';
partial_product_3(506) <= '0';
partial_product_3(507) <= '0';
partial_product_3(508) <= '0';
partial_product_3(509) <= '0';
partial_product_3(510) <= '0';
partial_product_3(511) <= '0';
partial_product_3(512) <= '0';
partial_product_4(0) <= '0';
partial_product_4(1) <= '0';
partial_product_4(2) <= '0';
partial_product_4(3) <= '0';
partial_product_4(4) <= '0';
partial_product_4(5) <= '0';
partial_product_4(6) <= '0';
partial_product_4(7) <= '0';
partial_product_4(8) <= '0';
partial_product_4(9) <= '0';
partial_product_4(10) <= '0';
partial_product_4(11) <= '0';
partial_product_4(12) <= '0';
partial_product_4(13) <= '0';
partial_product_4(14) <= '0';
partial_product_4(15) <= '0';
partial_product_4(16) <= '0';
partial_product_4(17) <= '0';
partial_product_4(18) <= '0';
partial_product_4(19) <= '0';
partial_product_4(20) <= '0';
partial_product_4(21) <= '0';
partial_product_4(22) <= '0';
partial_product_4(23) <= '0';
partial_product_4(24) <= '0';
partial_product_4(25) <= '0';
partial_product_4(26) <= '0';
partial_product_4(27) <= '0';
partial_product_4(28) <= '0';
partial_product_4(29) <= '0';
partial_product_4(30) <= '0';
partial_product_4(31) <= '0';
partial_product_4(32) <= '0';
partial_product_4(33) <= '0';
partial_product_4(34) <= '0';
partial_product_4(35) <= '0';
partial_product_4(36) <= '0';
partial_product_4(37) <= '0';
partial_product_4(38) <= '0';
partial_product_4(39) <= '0';
partial_product_4(40) <= '0';
partial_product_4(41) <= '0';
partial_product_4(42) <= '0';
partial_product_4(43) <= '0';
partial_product_4(44) <= '0';
partial_product_4(45) <= '0';
partial_product_4(46) <= '0';
partial_product_4(47) <= '0';
partial_product_4(48) <= temp_mult_2(48);
partial_product_4(49) <= temp_mult_2(49);
partial_product_4(50) <= temp_mult_2(50);
partial_product_4(51) <= temp_mult_2(51);
partial_product_4(52) <= temp_mult_2(52);
partial_product_4(53) <= temp_mult_2(53);
partial_product_4(54) <= temp_mult_2(54);
partial_product_4(55) <= temp_mult_2(55);
partial_product_4(56) <= temp_mult_2(56);
partial_product_4(57) <= temp_mult_2(57);
partial_product_4(58) <= temp_mult_2(58);
partial_product_4(59) <= temp_mult_2(59);
partial_product_4(60) <= temp_mult_2(60);
partial_product_4(61) <= temp_mult_2(61);
partial_product_4(62) <= temp_mult_2(62);
partial_product_4(63) <= temp_mult_2(63);
partial_product_4(64) <= temp_mult_2(64);
partial_product_4(65) <= temp_mult_2(65);
partial_product_4(66) <= temp_mult_2(66);
partial_product_4(67) <= temp_mult_2(67);
partial_product_4(68) <= temp_mult_2(68);
partial_product_4(69) <= temp_mult_2(69);
partial_product_4(70) <= temp_mult_2(70);
partial_product_4(71) <= temp_mult_2(71);
partial_product_4(72) <= temp_mult_2(72);
partial_product_4(73) <= temp_mult_2(73);
partial_product_4(74) <= temp_mult_2(74);
partial_product_4(75) <= temp_mult_2(75);
partial_product_4(76) <= temp_mult_2(76);
partial_product_4(77) <= temp_mult_2(77);
partial_product_4(78) <= temp_mult_2(78);
partial_product_4(79) <= temp_mult_2(79);
partial_product_4(80) <= temp_mult_2(80);
partial_product_4(81) <= temp_mult_2(81);
partial_product_4(82) <= temp_mult_2(82);
partial_product_4(83) <= temp_mult_2(83);
partial_product_4(84) <= temp_mult_2(84);
partial_product_4(85) <= temp_mult_2(85);
partial_product_4(86) <= temp_mult_2(86);
partial_product_4(87) <= temp_mult_2(87);
partial_product_4(88) <= temp_mult_2(88);
partial_product_4(89) <= temp_mult_8(89);
partial_product_4(90) <= temp_mult_8(90);
partial_product_4(91) <= temp_mult_8(91);
partial_product_4(92) <= temp_mult_8(92);
partial_product_4(93) <= temp_mult_8(93);
partial_product_4(94) <= temp_mult_8(94);
partial_product_4(95) <= temp_mult_8(95);
partial_product_4(96) <= temp_mult_8(96);
partial_product_4(97) <= temp_mult_8(97);
partial_product_4(98) <= temp_mult_8(98);
partial_product_4(99) <= temp_mult_8(99);
partial_product_4(100) <= temp_mult_8(100);
partial_product_4(101) <= temp_mult_8(101);
partial_product_4(102) <= temp_mult_8(102);
partial_product_4(103) <= temp_mult_8(103);
partial_product_4(104) <= temp_mult_8(104);
partial_product_4(105) <= temp_mult_8(105);
partial_product_4(106) <= temp_mult_8(106);
partial_product_4(107) <= temp_mult_8(107);
partial_product_4(108) <= temp_mult_8(108);
partial_product_4(109) <= temp_mult_8(109);
partial_product_4(110) <= temp_mult_8(110);
partial_product_4(111) <= temp_mult_8(111);
partial_product_4(112) <= temp_mult_8(112);
partial_product_4(113) <= temp_mult_8(113);
partial_product_4(114) <= temp_mult_8(114);
partial_product_4(115) <= temp_mult_8(115);
partial_product_4(116) <= temp_mult_8(116);
partial_product_4(117) <= temp_mult_8(117);
partial_product_4(118) <= temp_mult_8(118);
partial_product_4(119) <= temp_mult_8(119);
partial_product_4(120) <= temp_mult_8(120);
partial_product_4(121) <= temp_mult_8(121);
partial_product_4(122) <= temp_mult_8(122);
partial_product_4(123) <= temp_mult_8(123);
partial_product_4(124) <= temp_mult_8(124);
partial_product_4(125) <= temp_mult_8(125);
partial_product_4(126) <= temp_mult_8(126);
partial_product_4(127) <= temp_mult_8(127);
partial_product_4(128) <= temp_mult_8(128);
partial_product_4(129) <= temp_mult_8(129);
partial_product_4(130) <= temp_mult_14(130);
partial_product_4(131) <= temp_mult_14(131);
partial_product_4(132) <= temp_mult_14(132);
partial_product_4(133) <= temp_mult_14(133);
partial_product_4(134) <= temp_mult_14(134);
partial_product_4(135) <= temp_mult_14(135);
partial_product_4(136) <= temp_mult_14(136);
partial_product_4(137) <= temp_mult_14(137);
partial_product_4(138) <= temp_mult_14(138);
partial_product_4(139) <= temp_mult_14(139);
partial_product_4(140) <= temp_mult_14(140);
partial_product_4(141) <= temp_mult_14(141);
partial_product_4(142) <= temp_mult_14(142);
partial_product_4(143) <= temp_mult_14(143);
partial_product_4(144) <= temp_mult_14(144);
partial_product_4(145) <= temp_mult_14(145);
partial_product_4(146) <= temp_mult_14(146);
partial_product_4(147) <= temp_mult_14(147);
partial_product_4(148) <= temp_mult_14(148);
partial_product_4(149) <= temp_mult_14(149);
partial_product_4(150) <= temp_mult_14(150);
partial_product_4(151) <= temp_mult_14(151);
partial_product_4(152) <= temp_mult_14(152);
partial_product_4(153) <= temp_mult_14(153);
partial_product_4(154) <= temp_mult_14(154);
partial_product_4(155) <= temp_mult_14(155);
partial_product_4(156) <= temp_mult_14(156);
partial_product_4(157) <= temp_mult_14(157);
partial_product_4(158) <= temp_mult_14(158);
partial_product_4(159) <= temp_mult_14(159);
partial_product_4(160) <= temp_mult_14(160);
partial_product_4(161) <= temp_mult_14(161);
partial_product_4(162) <= temp_mult_14(162);
partial_product_4(163) <= temp_mult_14(163);
partial_product_4(164) <= temp_mult_14(164);
partial_product_4(165) <= temp_mult_14(165);
partial_product_4(166) <= temp_mult_14(166);
partial_product_4(167) <= temp_mult_14(167);
partial_product_4(168) <= temp_mult_14(168);
partial_product_4(169) <= temp_mult_14(169);
partial_product_4(170) <= temp_mult_14(170);
partial_product_4(171) <= temp_mult_43(171);
partial_product_4(172) <= temp_mult_43(172);
partial_product_4(173) <= temp_mult_43(173);
partial_product_4(174) <= temp_mult_43(174);
partial_product_4(175) <= temp_mult_43(175);
partial_product_4(176) <= temp_mult_43(176);
partial_product_4(177) <= temp_mult_43(177);
partial_product_4(178) <= temp_mult_43(178);
partial_product_4(179) <= temp_mult_43(179);
partial_product_4(180) <= temp_mult_43(180);
partial_product_4(181) <= temp_mult_43(181);
partial_product_4(182) <= temp_mult_43(182);
partial_product_4(183) <= temp_mult_43(183);
partial_product_4(184) <= temp_mult_43(184);
partial_product_4(185) <= temp_mult_43(185);
partial_product_4(186) <= temp_mult_43(186);
partial_product_4(187) <= temp_mult_43(187);
partial_product_4(188) <= temp_mult_43(188);
partial_product_4(189) <= temp_mult_43(189);
partial_product_4(190) <= temp_mult_43(190);
partial_product_4(191) <= temp_mult_43(191);
partial_product_4(192) <= temp_mult_43(192);
partial_product_4(193) <= temp_mult_43(193);
partial_product_4(194) <= temp_mult_43(194);
partial_product_4(195) <= temp_mult_43(195);
partial_product_4(196) <= temp_mult_43(196);
partial_product_4(197) <= temp_mult_43(197);
partial_product_4(198) <= temp_mult_43(198);
partial_product_4(199) <= temp_mult_43(199);
partial_product_4(200) <= temp_mult_43(200);
partial_product_4(201) <= temp_mult_43(201);
partial_product_4(202) <= temp_mult_43(202);
partial_product_4(203) <= temp_mult_43(203);
partial_product_4(204) <= temp_mult_43(204);
partial_product_4(205) <= temp_mult_43(205);
partial_product_4(206) <= temp_mult_43(206);
partial_product_4(207) <= temp_mult_43(207);
partial_product_4(208) <= temp_mult_43(208);
partial_product_4(209) <= temp_mult_43(209);
partial_product_4(210) <= temp_mult_43(210);
partial_product_4(211) <= temp_mult_43(211);
partial_product_4(212) <= temp_mult_52(212);
partial_product_4(213) <= temp_mult_52(213);
partial_product_4(214) <= temp_mult_52(214);
partial_product_4(215) <= temp_mult_52(215);
partial_product_4(216) <= temp_mult_52(216);
partial_product_4(217) <= temp_mult_52(217);
partial_product_4(218) <= temp_mult_52(218);
partial_product_4(219) <= temp_mult_52(219);
partial_product_4(220) <= temp_mult_52(220);
partial_product_4(221) <= temp_mult_52(221);
partial_product_4(222) <= temp_mult_52(222);
partial_product_4(223) <= temp_mult_52(223);
partial_product_4(224) <= temp_mult_52(224);
partial_product_4(225) <= temp_mult_52(225);
partial_product_4(226) <= temp_mult_52(226);
partial_product_4(227) <= temp_mult_52(227);
partial_product_4(228) <= temp_mult_52(228);
partial_product_4(229) <= temp_mult_52(229);
partial_product_4(230) <= temp_mult_52(230);
partial_product_4(231) <= temp_mult_52(231);
partial_product_4(232) <= temp_mult_52(232);
partial_product_4(233) <= temp_mult_52(233);
partial_product_4(234) <= temp_mult_52(234);
partial_product_4(235) <= temp_mult_52(235);
partial_product_4(236) <= temp_mult_52(236);
partial_product_4(237) <= temp_mult_52(237);
partial_product_4(238) <= temp_mult_52(238);
partial_product_4(239) <= temp_mult_52(239);
partial_product_4(240) <= temp_mult_52(240);
partial_product_4(241) <= temp_mult_52(241);
partial_product_4(242) <= temp_mult_52(242);
partial_product_4(243) <= temp_mult_52(243);
partial_product_4(244) <= temp_mult_52(244);
partial_product_4(245) <= temp_mult_52(245);
partial_product_4(246) <= temp_mult_52(246);
partial_product_4(247) <= temp_mult_52(247);
partial_product_4(248) <= temp_mult_52(248);
partial_product_4(249) <= temp_mult_52(249);
partial_product_4(250) <= temp_mult_52(250);
partial_product_4(251) <= temp_mult_52(251);
partial_product_4(252) <= temp_mult_52(252);
partial_product_4(253) <= temp_mult_61(253);
partial_product_4(254) <= temp_mult_61(254);
partial_product_4(255) <= temp_mult_61(255);
partial_product_4(256) <= temp_mult_61(256);
partial_product_4(257) <= temp_mult_61(257);
partial_product_4(258) <= temp_mult_61(258);
partial_product_4(259) <= temp_mult_61(259);
partial_product_4(260) <= temp_mult_61(260);
partial_product_4(261) <= temp_mult_61(261);
partial_product_4(262) <= temp_mult_61(262);
partial_product_4(263) <= temp_mult_61(263);
partial_product_4(264) <= temp_mult_61(264);
partial_product_4(265) <= temp_mult_61(265);
partial_product_4(266) <= temp_mult_61(266);
partial_product_4(267) <= temp_mult_61(267);
partial_product_4(268) <= temp_mult_61(268);
partial_product_4(269) <= temp_mult_61(269);
partial_product_4(270) <= temp_mult_61(270);
partial_product_4(271) <= temp_mult_61(271);
partial_product_4(272) <= temp_mult_61(272);
partial_product_4(273) <= temp_mult_61(273);
partial_product_4(274) <= temp_mult_61(274);
partial_product_4(275) <= temp_mult_61(275);
partial_product_4(276) <= temp_mult_61(276);
partial_product_4(277) <= temp_mult_61(277);
partial_product_4(278) <= temp_mult_61(278);
partial_product_4(279) <= temp_mult_61(279);
partial_product_4(280) <= temp_mult_61(280);
partial_product_4(281) <= temp_mult_61(281);
partial_product_4(282) <= temp_mult_61(282);
partial_product_4(283) <= temp_mult_61(283);
partial_product_4(284) <= temp_mult_61(284);
partial_product_4(285) <= temp_mult_61(285);
partial_product_4(286) <= temp_mult_61(286);
partial_product_4(287) <= temp_mult_61(287);
partial_product_4(288) <= temp_mult_61(288);
partial_product_4(289) <= temp_mult_61(289);
partial_product_4(290) <= temp_mult_61(290);
partial_product_4(291) <= temp_mult_61(291);
partial_product_4(292) <= temp_mult_61(292);
partial_product_4(293) <= temp_mult_61(293);
partial_product_4(294) <= temp_mult_70(294);
partial_product_4(295) <= temp_mult_70(295);
partial_product_4(296) <= temp_mult_70(296);
partial_product_4(297) <= temp_mult_70(297);
partial_product_4(298) <= temp_mult_70(298);
partial_product_4(299) <= temp_mult_70(299);
partial_product_4(300) <= temp_mult_70(300);
partial_product_4(301) <= temp_mult_70(301);
partial_product_4(302) <= temp_mult_70(302);
partial_product_4(303) <= temp_mult_70(303);
partial_product_4(304) <= temp_mult_70(304);
partial_product_4(305) <= temp_mult_70(305);
partial_product_4(306) <= temp_mult_70(306);
partial_product_4(307) <= temp_mult_70(307);
partial_product_4(308) <= temp_mult_70(308);
partial_product_4(309) <= temp_mult_70(309);
partial_product_4(310) <= temp_mult_70(310);
partial_product_4(311) <= temp_mult_70(311);
partial_product_4(312) <= temp_mult_70(312);
partial_product_4(313) <= temp_mult_70(313);
partial_product_4(314) <= temp_mult_70(314);
partial_product_4(315) <= temp_mult_70(315);
partial_product_4(316) <= temp_mult_70(316);
partial_product_4(317) <= temp_mult_70(317);
partial_product_4(318) <= temp_mult_70(318);
partial_product_4(319) <= temp_mult_70(319);
partial_product_4(320) <= temp_mult_70(320);
partial_product_4(321) <= temp_mult_70(321);
partial_product_4(322) <= temp_mult_70(322);
partial_product_4(323) <= temp_mult_70(323);
partial_product_4(324) <= temp_mult_70(324);
partial_product_4(325) <= temp_mult_70(325);
partial_product_4(326) <= temp_mult_70(326);
partial_product_4(327) <= temp_mult_70(327);
partial_product_4(328) <= temp_mult_70(328);
partial_product_4(329) <= temp_mult_70(329);
partial_product_4(330) <= temp_mult_70(330);
partial_product_4(331) <= temp_mult_70(331);
partial_product_4(332) <= temp_mult_70(332);
partial_product_4(333) <= temp_mult_70(333);
partial_product_4(334) <= temp_mult_70(334);
partial_product_4(335) <= temp_mult_79(335);
partial_product_4(336) <= temp_mult_79(336);
partial_product_4(337) <= temp_mult_79(337);
partial_product_4(338) <= temp_mult_79(338);
partial_product_4(339) <= temp_mult_79(339);
partial_product_4(340) <= temp_mult_79(340);
partial_product_4(341) <= temp_mult_79(341);
partial_product_4(342) <= temp_mult_79(342);
partial_product_4(343) <= temp_mult_79(343);
partial_product_4(344) <= temp_mult_79(344);
partial_product_4(345) <= temp_mult_79(345);
partial_product_4(346) <= temp_mult_79(346);
partial_product_4(347) <= temp_mult_79(347);
partial_product_4(348) <= temp_mult_79(348);
partial_product_4(349) <= temp_mult_79(349);
partial_product_4(350) <= temp_mult_79(350);
partial_product_4(351) <= temp_mult_79(351);
partial_product_4(352) <= temp_mult_79(352);
partial_product_4(353) <= temp_mult_79(353);
partial_product_4(354) <= temp_mult_79(354);
partial_product_4(355) <= temp_mult_79(355);
partial_product_4(356) <= temp_mult_79(356);
partial_product_4(357) <= temp_mult_79(357);
partial_product_4(358) <= temp_mult_79(358);
partial_product_4(359) <= temp_mult_79(359);
partial_product_4(360) <= temp_mult_79(360);
partial_product_4(361) <= temp_mult_79(361);
partial_product_4(362) <= temp_mult_79(362);
partial_product_4(363) <= temp_mult_79(363);
partial_product_4(364) <= temp_mult_79(364);
partial_product_4(365) <= temp_mult_79(365);
partial_product_4(366) <= temp_mult_79(366);
partial_product_4(367) <= temp_mult_79(367);
partial_product_4(368) <= temp_mult_79(368);
partial_product_4(369) <= temp_mult_79(369);
partial_product_4(370) <= temp_mult_79(370);
partial_product_4(371) <= temp_mult_79(371);
partial_product_4(372) <= temp_mult_79(372);
partial_product_4(373) <= temp_mult_79(373);
partial_product_4(374) <= temp_mult_79(374);
partial_product_4(375) <= temp_mult_79(375);
partial_product_4(376) <= '0';
partial_product_4(377) <= '0';
partial_product_4(378) <= '0';
partial_product_4(379) <= temp_mult_138(379);
partial_product_4(380) <= temp_mult_138(380);
partial_product_4(381) <= temp_mult_138(381);
partial_product_4(382) <= temp_mult_138(382);
partial_product_4(383) <= temp_mult_138(383);
partial_product_4(384) <= temp_mult_138(384);
partial_product_4(385) <= temp_mult_138(385);
partial_product_4(386) <= temp_mult_138(386);
partial_product_4(387) <= temp_mult_138(387);
partial_product_4(388) <= temp_mult_138(388);
partial_product_4(389) <= temp_mult_138(389);
partial_product_4(390) <= temp_mult_138(390);
partial_product_4(391) <= temp_mult_138(391);
partial_product_4(392) <= temp_mult_138(392);
partial_product_4(393) <= temp_mult_138(393);
partial_product_4(394) <= temp_mult_138(394);
partial_product_4(395) <= temp_mult_138(395);
partial_product_4(396) <= temp_mult_138(396);
partial_product_4(397) <= temp_mult_138(397);
partial_product_4(398) <= temp_mult_138(398);
partial_product_4(399) <= temp_mult_138(399);
partial_product_4(400) <= temp_mult_138(400);
partial_product_4(401) <= temp_mult_138(401);
partial_product_4(402) <= temp_mult_138(402);
partial_product_4(403) <= temp_mult_138(403);
partial_product_4(404) <= temp_mult_138(404);
partial_product_4(405) <= temp_mult_138(405);
partial_product_4(406) <= temp_mult_138(406);
partial_product_4(407) <= temp_mult_138(407);
partial_product_4(408) <= temp_mult_138(408);
partial_product_4(409) <= temp_mult_138(409);
partial_product_4(410) <= temp_mult_138(410);
partial_product_4(411) <= temp_mult_138(411);
partial_product_4(412) <= temp_mult_138(412);
partial_product_4(413) <= temp_mult_138(413);
partial_product_4(414) <= temp_mult_138(414);
partial_product_4(415) <= temp_mult_138(415);
partial_product_4(416) <= temp_mult_138(416);
partial_product_4(417) <= temp_mult_138(417);
partial_product_4(418) <= temp_mult_138(418);
partial_product_4(419) <= temp_mult_138(419);
partial_product_4(420) <= temp_mult_144(420);
partial_product_4(421) <= temp_mult_144(421);
partial_product_4(422) <= temp_mult_144(422);
partial_product_4(423) <= temp_mult_144(423);
partial_product_4(424) <= temp_mult_144(424);
partial_product_4(425) <= temp_mult_144(425);
partial_product_4(426) <= temp_mult_144(426);
partial_product_4(427) <= temp_mult_144(427);
partial_product_4(428) <= temp_mult_144(428);
partial_product_4(429) <= temp_mult_144(429);
partial_product_4(430) <= temp_mult_144(430);
partial_product_4(431) <= temp_mult_144(431);
partial_product_4(432) <= temp_mult_144(432);
partial_product_4(433) <= temp_mult_144(433);
partial_product_4(434) <= temp_mult_144(434);
partial_product_4(435) <= temp_mult_144(435);
partial_product_4(436) <= temp_mult_144(436);
partial_product_4(437) <= temp_mult_144(437);
partial_product_4(438) <= temp_mult_144(438);
partial_product_4(439) <= temp_mult_144(439);
partial_product_4(440) <= temp_mult_144(440);
partial_product_4(441) <= temp_mult_144(441);
partial_product_4(442) <= temp_mult_144(442);
partial_product_4(443) <= temp_mult_144(443);
partial_product_4(444) <= temp_mult_144(444);
partial_product_4(445) <= temp_mult_144(445);
partial_product_4(446) <= temp_mult_144(446);
partial_product_4(447) <= temp_mult_144(447);
partial_product_4(448) <= temp_mult_144(448);
partial_product_4(449) <= temp_mult_144(449);
partial_product_4(450) <= temp_mult_144(450);
partial_product_4(451) <= temp_mult_144(451);
partial_product_4(452) <= temp_mult_144(452);
partial_product_4(453) <= temp_mult_144(453);
partial_product_4(454) <= temp_mult_144(454);
partial_product_4(455) <= temp_mult_144(455);
partial_product_4(456) <= temp_mult_144(456);
partial_product_4(457) <= temp_mult_144(457);
partial_product_4(458) <= temp_mult_144(458);
partial_product_4(459) <= temp_mult_144(459);
partial_product_4(460) <= temp_mult_144(460);
partial_product_4(461) <= '0';
partial_product_4(462) <= '0';
partial_product_4(463) <= '0';
partial_product_4(464) <= '0';
partial_product_4(465) <= '0';
partial_product_4(466) <= '0';
partial_product_4(467) <= '0';
partial_product_4(468) <= '0';
partial_product_4(469) <= '0';
partial_product_4(470) <= '0';
partial_product_4(471) <= '0';
partial_product_4(472) <= '0';
partial_product_4(473) <= '0';
partial_product_4(474) <= '0';
partial_product_4(475) <= '0';
partial_product_4(476) <= '0';
partial_product_4(477) <= '0';
partial_product_4(478) <= '0';
partial_product_4(479) <= '0';
partial_product_4(480) <= '0';
partial_product_4(481) <= '0';
partial_product_4(482) <= '0';
partial_product_4(483) <= '0';
partial_product_4(484) <= '0';
partial_product_4(485) <= '0';
partial_product_4(486) <= '0';
partial_product_4(487) <= '0';
partial_product_4(488) <= '0';
partial_product_4(489) <= '0';
partial_product_4(490) <= '0';
partial_product_4(491) <= '0';
partial_product_4(492) <= '0';
partial_product_4(493) <= '0';
partial_product_4(494) <= '0';
partial_product_4(495) <= '0';
partial_product_4(496) <= '0';
partial_product_4(497) <= '0';
partial_product_4(498) <= '0';
partial_product_4(499) <= '0';
partial_product_4(500) <= '0';
partial_product_4(501) <= '0';
partial_product_4(502) <= '0';
partial_product_4(503) <= '0';
partial_product_4(504) <= '0';
partial_product_4(505) <= '0';
partial_product_4(506) <= '0';
partial_product_4(507) <= '0';
partial_product_4(508) <= '0';
partial_product_4(509) <= '0';
partial_product_4(510) <= '0';
partial_product_4(511) <= '0';
partial_product_4(512) <= '0';
partial_product_5(0) <= '0';
partial_product_5(1) <= '0';
partial_product_5(2) <= '0';
partial_product_5(3) <= '0';
partial_product_5(4) <= '0';
partial_product_5(5) <= '0';
partial_product_5(6) <= '0';
partial_product_5(7) <= '0';
partial_product_5(8) <= '0';
partial_product_5(9) <= '0';
partial_product_5(10) <= '0';
partial_product_5(11) <= '0';
partial_product_5(12) <= '0';
partial_product_5(13) <= '0';
partial_product_5(14) <= '0';
partial_product_5(15) <= '0';
partial_product_5(16) <= '0';
partial_product_5(17) <= '0';
partial_product_5(18) <= '0';
partial_product_5(19) <= '0';
partial_product_5(20) <= '0';
partial_product_5(21) <= '0';
partial_product_5(22) <= '0';
partial_product_5(23) <= '0';
partial_product_5(24) <= '0';
partial_product_5(25) <= '0';
partial_product_5(26) <= '0';
partial_product_5(27) <= '0';
partial_product_5(28) <= '0';
partial_product_5(29) <= '0';
partial_product_5(30) <= '0';
partial_product_5(31) <= '0';
partial_product_5(32) <= '0';
partial_product_5(33) <= '0';
partial_product_5(34) <= '0';
partial_product_5(35) <= '0';
partial_product_5(36) <= '0';
partial_product_5(37) <= '0';
partial_product_5(38) <= '0';
partial_product_5(39) <= '0';
partial_product_5(40) <= '0';
partial_product_5(41) <= '0';
partial_product_5(42) <= '0';
partial_product_5(43) <= '0';
partial_product_5(44) <= '0';
partial_product_5(45) <= '0';
partial_product_5(46) <= '0';
partial_product_5(47) <= '0';
partial_product_5(48) <= '0';
partial_product_5(49) <= '0';
partial_product_5(50) <= '0';
partial_product_5(51) <= temp_mult_15(51);
partial_product_5(52) <= temp_mult_15(52);
partial_product_5(53) <= temp_mult_15(53);
partial_product_5(54) <= temp_mult_15(54);
partial_product_5(55) <= temp_mult_15(55);
partial_product_5(56) <= temp_mult_15(56);
partial_product_5(57) <= temp_mult_15(57);
partial_product_5(58) <= temp_mult_15(58);
partial_product_5(59) <= temp_mult_15(59);
partial_product_5(60) <= temp_mult_15(60);
partial_product_5(61) <= temp_mult_15(61);
partial_product_5(62) <= temp_mult_15(62);
partial_product_5(63) <= temp_mult_15(63);
partial_product_5(64) <= temp_mult_15(64);
partial_product_5(65) <= temp_mult_15(65);
partial_product_5(66) <= temp_mult_15(66);
partial_product_5(67) <= temp_mult_15(67);
partial_product_5(68) <= temp_mult_15(68);
partial_product_5(69) <= temp_mult_15(69);
partial_product_5(70) <= temp_mult_15(70);
partial_product_5(71) <= temp_mult_15(71);
partial_product_5(72) <= temp_mult_15(72);
partial_product_5(73) <= temp_mult_15(73);
partial_product_5(74) <= temp_mult_15(74);
partial_product_5(75) <= temp_mult_15(75);
partial_product_5(76) <= temp_mult_15(76);
partial_product_5(77) <= temp_mult_15(77);
partial_product_5(78) <= temp_mult_15(78);
partial_product_5(79) <= temp_mult_15(79);
partial_product_5(80) <= temp_mult_15(80);
partial_product_5(81) <= temp_mult_15(81);
partial_product_5(82) <= temp_mult_15(82);
partial_product_5(83) <= temp_mult_15(83);
partial_product_5(84) <= temp_mult_15(84);
partial_product_5(85) <= temp_mult_15(85);
partial_product_5(86) <= temp_mult_15(86);
partial_product_5(87) <= temp_mult_15(87);
partial_product_5(88) <= temp_mult_15(88);
partial_product_5(89) <= temp_mult_15(89);
partial_product_5(90) <= temp_mult_15(90);
partial_product_5(91) <= temp_mult_15(91);
partial_product_5(92) <= temp_mult_21(92);
partial_product_5(93) <= temp_mult_21(93);
partial_product_5(94) <= temp_mult_21(94);
partial_product_5(95) <= temp_mult_21(95);
partial_product_5(96) <= temp_mult_21(96);
partial_product_5(97) <= temp_mult_21(97);
partial_product_5(98) <= temp_mult_21(98);
partial_product_5(99) <= temp_mult_21(99);
partial_product_5(100) <= temp_mult_21(100);
partial_product_5(101) <= temp_mult_21(101);
partial_product_5(102) <= temp_mult_21(102);
partial_product_5(103) <= temp_mult_21(103);
partial_product_5(104) <= temp_mult_21(104);
partial_product_5(105) <= temp_mult_21(105);
partial_product_5(106) <= temp_mult_21(106);
partial_product_5(107) <= temp_mult_21(107);
partial_product_5(108) <= temp_mult_21(108);
partial_product_5(109) <= temp_mult_21(109);
partial_product_5(110) <= temp_mult_21(110);
partial_product_5(111) <= temp_mult_21(111);
partial_product_5(112) <= temp_mult_21(112);
partial_product_5(113) <= temp_mult_21(113);
partial_product_5(114) <= temp_mult_21(114);
partial_product_5(115) <= temp_mult_21(115);
partial_product_5(116) <= temp_mult_21(116);
partial_product_5(117) <= temp_mult_21(117);
partial_product_5(118) <= temp_mult_21(118);
partial_product_5(119) <= temp_mult_21(119);
partial_product_5(120) <= temp_mult_21(120);
partial_product_5(121) <= temp_mult_21(121);
partial_product_5(122) <= temp_mult_21(122);
partial_product_5(123) <= temp_mult_21(123);
partial_product_5(124) <= temp_mult_21(124);
partial_product_5(125) <= temp_mult_21(125);
partial_product_5(126) <= temp_mult_21(126);
partial_product_5(127) <= temp_mult_21(127);
partial_product_5(128) <= temp_mult_21(128);
partial_product_5(129) <= temp_mult_21(129);
partial_product_5(130) <= temp_mult_21(130);
partial_product_5(131) <= temp_mult_21(131);
partial_product_5(132) <= temp_mult_21(132);
partial_product_5(133) <= temp_mult_27(133);
partial_product_5(134) <= temp_mult_27(134);
partial_product_5(135) <= temp_mult_27(135);
partial_product_5(136) <= temp_mult_27(136);
partial_product_5(137) <= temp_mult_27(137);
partial_product_5(138) <= temp_mult_27(138);
partial_product_5(139) <= temp_mult_27(139);
partial_product_5(140) <= temp_mult_27(140);
partial_product_5(141) <= temp_mult_27(141);
partial_product_5(142) <= temp_mult_27(142);
partial_product_5(143) <= temp_mult_27(143);
partial_product_5(144) <= temp_mult_27(144);
partial_product_5(145) <= temp_mult_27(145);
partial_product_5(146) <= temp_mult_27(146);
partial_product_5(147) <= temp_mult_27(147);
partial_product_5(148) <= temp_mult_27(148);
partial_product_5(149) <= temp_mult_27(149);
partial_product_5(150) <= temp_mult_27(150);
partial_product_5(151) <= temp_mult_27(151);
partial_product_5(152) <= temp_mult_27(152);
partial_product_5(153) <= temp_mult_27(153);
partial_product_5(154) <= temp_mult_27(154);
partial_product_5(155) <= temp_mult_27(155);
partial_product_5(156) <= temp_mult_27(156);
partial_product_5(157) <= temp_mult_27(157);
partial_product_5(158) <= temp_mult_27(158);
partial_product_5(159) <= temp_mult_27(159);
partial_product_5(160) <= temp_mult_27(160);
partial_product_5(161) <= temp_mult_27(161);
partial_product_5(162) <= temp_mult_27(162);
partial_product_5(163) <= temp_mult_27(163);
partial_product_5(164) <= temp_mult_27(164);
partial_product_5(165) <= temp_mult_27(165);
partial_product_5(166) <= temp_mult_27(166);
partial_product_5(167) <= temp_mult_27(167);
partial_product_5(168) <= temp_mult_27(168);
partial_product_5(169) <= temp_mult_27(169);
partial_product_5(170) <= temp_mult_27(170);
partial_product_5(171) <= temp_mult_27(171);
partial_product_5(172) <= temp_mult_27(172);
partial_product_5(173) <= temp_mult_27(173);
partial_product_5(174) <= temp_mult_33(174);
partial_product_5(175) <= temp_mult_33(175);
partial_product_5(176) <= temp_mult_33(176);
partial_product_5(177) <= temp_mult_33(177);
partial_product_5(178) <= temp_mult_33(178);
partial_product_5(179) <= temp_mult_33(179);
partial_product_5(180) <= temp_mult_33(180);
partial_product_5(181) <= temp_mult_33(181);
partial_product_5(182) <= temp_mult_33(182);
partial_product_5(183) <= temp_mult_33(183);
partial_product_5(184) <= temp_mult_33(184);
partial_product_5(185) <= temp_mult_33(185);
partial_product_5(186) <= temp_mult_33(186);
partial_product_5(187) <= temp_mult_33(187);
partial_product_5(188) <= temp_mult_33(188);
partial_product_5(189) <= temp_mult_33(189);
partial_product_5(190) <= temp_mult_33(190);
partial_product_5(191) <= temp_mult_33(191);
partial_product_5(192) <= temp_mult_33(192);
partial_product_5(193) <= temp_mult_33(193);
partial_product_5(194) <= temp_mult_33(194);
partial_product_5(195) <= temp_mult_33(195);
partial_product_5(196) <= temp_mult_33(196);
partial_product_5(197) <= temp_mult_33(197);
partial_product_5(198) <= temp_mult_33(198);
partial_product_5(199) <= temp_mult_33(199);
partial_product_5(200) <= temp_mult_33(200);
partial_product_5(201) <= temp_mult_33(201);
partial_product_5(202) <= temp_mult_33(202);
partial_product_5(203) <= temp_mult_33(203);
partial_product_5(204) <= temp_mult_33(204);
partial_product_5(205) <= temp_mult_33(205);
partial_product_5(206) <= temp_mult_33(206);
partial_product_5(207) <= temp_mult_33(207);
partial_product_5(208) <= temp_mult_33(208);
partial_product_5(209) <= temp_mult_33(209);
partial_product_5(210) <= temp_mult_33(210);
partial_product_5(211) <= temp_mult_33(211);
partial_product_5(212) <= temp_mult_33(212);
partial_product_5(213) <= temp_mult_33(213);
partial_product_5(214) <= temp_mult_33(214);
partial_product_5(215) <= temp_mult_39(215);
partial_product_5(216) <= temp_mult_39(216);
partial_product_5(217) <= temp_mult_39(217);
partial_product_5(218) <= temp_mult_39(218);
partial_product_5(219) <= temp_mult_39(219);
partial_product_5(220) <= temp_mult_39(220);
partial_product_5(221) <= temp_mult_39(221);
partial_product_5(222) <= temp_mult_39(222);
partial_product_5(223) <= temp_mult_39(223);
partial_product_5(224) <= temp_mult_39(224);
partial_product_5(225) <= temp_mult_39(225);
partial_product_5(226) <= temp_mult_39(226);
partial_product_5(227) <= temp_mult_39(227);
partial_product_5(228) <= temp_mult_39(228);
partial_product_5(229) <= temp_mult_39(229);
partial_product_5(230) <= temp_mult_39(230);
partial_product_5(231) <= temp_mult_39(231);
partial_product_5(232) <= temp_mult_39(232);
partial_product_5(233) <= temp_mult_39(233);
partial_product_5(234) <= temp_mult_39(234);
partial_product_5(235) <= temp_mult_39(235);
partial_product_5(236) <= temp_mult_39(236);
partial_product_5(237) <= temp_mult_39(237);
partial_product_5(238) <= temp_mult_39(238);
partial_product_5(239) <= temp_mult_39(239);
partial_product_5(240) <= temp_mult_39(240);
partial_product_5(241) <= temp_mult_39(241);
partial_product_5(242) <= temp_mult_39(242);
partial_product_5(243) <= temp_mult_39(243);
partial_product_5(244) <= temp_mult_39(244);
partial_product_5(245) <= temp_mult_39(245);
partial_product_5(246) <= temp_mult_39(246);
partial_product_5(247) <= temp_mult_39(247);
partial_product_5(248) <= temp_mult_39(248);
partial_product_5(249) <= temp_mult_39(249);
partial_product_5(250) <= temp_mult_39(250);
partial_product_5(251) <= temp_mult_39(251);
partial_product_5(252) <= temp_mult_39(252);
partial_product_5(253) <= temp_mult_39(253);
partial_product_5(254) <= temp_mult_39(254);
partial_product_5(255) <= temp_mult_39(255);
partial_product_5(256) <= temp_mult_120(256);
partial_product_5(257) <= temp_mult_120(257);
partial_product_5(258) <= temp_mult_120(258);
partial_product_5(259) <= temp_mult_120(259);
partial_product_5(260) <= temp_mult_120(260);
partial_product_5(261) <= temp_mult_120(261);
partial_product_5(262) <= temp_mult_120(262);
partial_product_5(263) <= temp_mult_120(263);
partial_product_5(264) <= temp_mult_120(264);
partial_product_5(265) <= temp_mult_120(265);
partial_product_5(266) <= temp_mult_120(266);
partial_product_5(267) <= temp_mult_120(267);
partial_product_5(268) <= temp_mult_120(268);
partial_product_5(269) <= temp_mult_120(269);
partial_product_5(270) <= temp_mult_120(270);
partial_product_5(271) <= temp_mult_120(271);
partial_product_5(272) <= temp_mult_120(272);
partial_product_5(273) <= temp_mult_120(273);
partial_product_5(274) <= temp_mult_120(274);
partial_product_5(275) <= temp_mult_120(275);
partial_product_5(276) <= temp_mult_120(276);
partial_product_5(277) <= temp_mult_120(277);
partial_product_5(278) <= temp_mult_120(278);
partial_product_5(279) <= temp_mult_120(279);
partial_product_5(280) <= temp_mult_120(280);
partial_product_5(281) <= temp_mult_120(281);
partial_product_5(282) <= temp_mult_120(282);
partial_product_5(283) <= temp_mult_120(283);
partial_product_5(284) <= temp_mult_120(284);
partial_product_5(285) <= temp_mult_120(285);
partial_product_5(286) <= temp_mult_120(286);
partial_product_5(287) <= temp_mult_120(287);
partial_product_5(288) <= temp_mult_120(288);
partial_product_5(289) <= temp_mult_120(289);
partial_product_5(290) <= temp_mult_120(290);
partial_product_5(291) <= temp_mult_120(291);
partial_product_5(292) <= temp_mult_120(292);
partial_product_5(293) <= temp_mult_120(293);
partial_product_5(294) <= temp_mult_120(294);
partial_product_5(295) <= temp_mult_120(295);
partial_product_5(296) <= temp_mult_120(296);
partial_product_5(297) <= temp_mult_126(297);
partial_product_5(298) <= temp_mult_126(298);
partial_product_5(299) <= temp_mult_126(299);
partial_product_5(300) <= temp_mult_126(300);
partial_product_5(301) <= temp_mult_126(301);
partial_product_5(302) <= temp_mult_126(302);
partial_product_5(303) <= temp_mult_126(303);
partial_product_5(304) <= temp_mult_126(304);
partial_product_5(305) <= temp_mult_126(305);
partial_product_5(306) <= temp_mult_126(306);
partial_product_5(307) <= temp_mult_126(307);
partial_product_5(308) <= temp_mult_126(308);
partial_product_5(309) <= temp_mult_126(309);
partial_product_5(310) <= temp_mult_126(310);
partial_product_5(311) <= temp_mult_126(311);
partial_product_5(312) <= temp_mult_126(312);
partial_product_5(313) <= temp_mult_126(313);
partial_product_5(314) <= temp_mult_126(314);
partial_product_5(315) <= temp_mult_126(315);
partial_product_5(316) <= temp_mult_126(316);
partial_product_5(317) <= temp_mult_126(317);
partial_product_5(318) <= temp_mult_126(318);
partial_product_5(319) <= temp_mult_126(319);
partial_product_5(320) <= temp_mult_126(320);
partial_product_5(321) <= temp_mult_126(321);
partial_product_5(322) <= temp_mult_126(322);
partial_product_5(323) <= temp_mult_126(323);
partial_product_5(324) <= temp_mult_126(324);
partial_product_5(325) <= temp_mult_126(325);
partial_product_5(326) <= temp_mult_126(326);
partial_product_5(327) <= temp_mult_126(327);
partial_product_5(328) <= temp_mult_126(328);
partial_product_5(329) <= temp_mult_126(329);
partial_product_5(330) <= temp_mult_126(330);
partial_product_5(331) <= temp_mult_126(331);
partial_product_5(332) <= temp_mult_126(332);
partial_product_5(333) <= temp_mult_126(333);
partial_product_5(334) <= temp_mult_126(334);
partial_product_5(335) <= temp_mult_126(335);
partial_product_5(336) <= temp_mult_126(336);
partial_product_5(337) <= temp_mult_126(337);
partial_product_5(338) <= temp_mult_132(338);
partial_product_5(339) <= temp_mult_132(339);
partial_product_5(340) <= temp_mult_132(340);
partial_product_5(341) <= temp_mult_132(341);
partial_product_5(342) <= temp_mult_132(342);
partial_product_5(343) <= temp_mult_132(343);
partial_product_5(344) <= temp_mult_132(344);
partial_product_5(345) <= temp_mult_132(345);
partial_product_5(346) <= temp_mult_132(346);
partial_product_5(347) <= temp_mult_132(347);
partial_product_5(348) <= temp_mult_132(348);
partial_product_5(349) <= temp_mult_132(349);
partial_product_5(350) <= temp_mult_132(350);
partial_product_5(351) <= temp_mult_132(351);
partial_product_5(352) <= temp_mult_132(352);
partial_product_5(353) <= temp_mult_132(353);
partial_product_5(354) <= temp_mult_132(354);
partial_product_5(355) <= temp_mult_132(355);
partial_product_5(356) <= temp_mult_132(356);
partial_product_5(357) <= temp_mult_132(357);
partial_product_5(358) <= temp_mult_132(358);
partial_product_5(359) <= temp_mult_132(359);
partial_product_5(360) <= temp_mult_132(360);
partial_product_5(361) <= temp_mult_132(361);
partial_product_5(362) <= temp_mult_132(362);
partial_product_5(363) <= temp_mult_132(363);
partial_product_5(364) <= temp_mult_132(364);
partial_product_5(365) <= temp_mult_132(365);
partial_product_5(366) <= temp_mult_132(366);
partial_product_5(367) <= temp_mult_132(367);
partial_product_5(368) <= temp_mult_132(368);
partial_product_5(369) <= temp_mult_132(369);
partial_product_5(370) <= temp_mult_132(370);
partial_product_5(371) <= temp_mult_132(371);
partial_product_5(372) <= temp_mult_132(372);
partial_product_5(373) <= temp_mult_132(373);
partial_product_5(374) <= temp_mult_132(374);
partial_product_5(375) <= temp_mult_132(375);
partial_product_5(376) <= temp_mult_132(376);
partial_product_5(377) <= temp_mult_132(377);
partial_product_5(378) <= temp_mult_132(378);
partial_product_5(379) <= '0';
partial_product_5(380) <= '0';
partial_product_5(381) <= '0';
partial_product_5(382) <= temp_mult_151(382);
partial_product_5(383) <= temp_mult_151(383);
partial_product_5(384) <= temp_mult_151(384);
partial_product_5(385) <= temp_mult_151(385);
partial_product_5(386) <= temp_mult_151(386);
partial_product_5(387) <= temp_mult_151(387);
partial_product_5(388) <= temp_mult_151(388);
partial_product_5(389) <= temp_mult_151(389);
partial_product_5(390) <= temp_mult_151(390);
partial_product_5(391) <= temp_mult_151(391);
partial_product_5(392) <= temp_mult_151(392);
partial_product_5(393) <= temp_mult_151(393);
partial_product_5(394) <= temp_mult_151(394);
partial_product_5(395) <= temp_mult_151(395);
partial_product_5(396) <= temp_mult_151(396);
partial_product_5(397) <= temp_mult_151(397);
partial_product_5(398) <= temp_mult_151(398);
partial_product_5(399) <= temp_mult_151(399);
partial_product_5(400) <= temp_mult_151(400);
partial_product_5(401) <= temp_mult_151(401);
partial_product_5(402) <= temp_mult_151(402);
partial_product_5(403) <= temp_mult_151(403);
partial_product_5(404) <= temp_mult_151(404);
partial_product_5(405) <= temp_mult_151(405);
partial_product_5(406) <= temp_mult_151(406);
partial_product_5(407) <= temp_mult_151(407);
partial_product_5(408) <= temp_mult_151(408);
partial_product_5(409) <= temp_mult_151(409);
partial_product_5(410) <= temp_mult_151(410);
partial_product_5(411) <= temp_mult_151(411);
partial_product_5(412) <= temp_mult_151(412);
partial_product_5(413) <= temp_mult_151(413);
partial_product_5(414) <= temp_mult_151(414);
partial_product_5(415) <= temp_mult_151(415);
partial_product_5(416) <= temp_mult_151(416);
partial_product_5(417) <= temp_mult_151(417);
partial_product_5(418) <= temp_mult_151(418);
partial_product_5(419) <= temp_mult_151(419);
partial_product_5(420) <= temp_mult_151(420);
partial_product_5(421) <= temp_mult_151(421);
partial_product_5(422) <= temp_mult_151(422);
partial_product_5(423) <= temp_mult_157(423);
partial_product_5(424) <= temp_mult_157(424);
partial_product_5(425) <= temp_mult_157(425);
partial_product_5(426) <= temp_mult_157(426);
partial_product_5(427) <= temp_mult_157(427);
partial_product_5(428) <= temp_mult_157(428);
partial_product_5(429) <= temp_mult_157(429);
partial_product_5(430) <= temp_mult_157(430);
partial_product_5(431) <= temp_mult_157(431);
partial_product_5(432) <= temp_mult_157(432);
partial_product_5(433) <= temp_mult_157(433);
partial_product_5(434) <= temp_mult_157(434);
partial_product_5(435) <= temp_mult_157(435);
partial_product_5(436) <= temp_mult_157(436);
partial_product_5(437) <= temp_mult_157(437);
partial_product_5(438) <= temp_mult_157(438);
partial_product_5(439) <= temp_mult_157(439);
partial_product_5(440) <= temp_mult_157(440);
partial_product_5(441) <= temp_mult_157(441);
partial_product_5(442) <= temp_mult_157(442);
partial_product_5(443) <= temp_mult_157(443);
partial_product_5(444) <= temp_mult_157(444);
partial_product_5(445) <= temp_mult_157(445);
partial_product_5(446) <= temp_mult_157(446);
partial_product_5(447) <= temp_mult_157(447);
partial_product_5(448) <= temp_mult_157(448);
partial_product_5(449) <= temp_mult_157(449);
partial_product_5(450) <= temp_mult_157(450);
partial_product_5(451) <= temp_mult_157(451);
partial_product_5(452) <= temp_mult_157(452);
partial_product_5(453) <= temp_mult_157(453);
partial_product_5(454) <= temp_mult_157(454);
partial_product_5(455) <= temp_mult_157(455);
partial_product_5(456) <= temp_mult_157(456);
partial_product_5(457) <= temp_mult_157(457);
partial_product_5(458) <= temp_mult_157(458);
partial_product_5(459) <= temp_mult_157(459);
partial_product_5(460) <= temp_mult_157(460);
partial_product_5(461) <= temp_mult_157(461);
partial_product_5(462) <= temp_mult_157(462);
partial_product_5(463) <= temp_mult_157(463);
partial_product_5(464) <= '0';
partial_product_5(465) <= '0';
partial_product_5(466) <= '0';
partial_product_5(467) <= '0';
partial_product_5(468) <= '0';
partial_product_5(469) <= '0';
partial_product_5(470) <= '0';
partial_product_5(471) <= '0';
partial_product_5(472) <= '0';
partial_product_5(473) <= '0';
partial_product_5(474) <= '0';
partial_product_5(475) <= '0';
partial_product_5(476) <= '0';
partial_product_5(477) <= '0';
partial_product_5(478) <= '0';
partial_product_5(479) <= '0';
partial_product_5(480) <= '0';
partial_product_5(481) <= '0';
partial_product_5(482) <= '0';
partial_product_5(483) <= '0';
partial_product_5(484) <= '0';
partial_product_5(485) <= '0';
partial_product_5(486) <= '0';
partial_product_5(487) <= '0';
partial_product_5(488) <= '0';
partial_product_5(489) <= '0';
partial_product_5(490) <= '0';
partial_product_5(491) <= '0';
partial_product_5(492) <= '0';
partial_product_5(493) <= '0';
partial_product_5(494) <= '0';
partial_product_5(495) <= '0';
partial_product_5(496) <= '0';
partial_product_5(497) <= '0';
partial_product_5(498) <= '0';
partial_product_5(499) <= '0';
partial_product_5(500) <= '0';
partial_product_5(501) <= '0';
partial_product_5(502) <= '0';
partial_product_5(503) <= '0';
partial_product_5(504) <= '0';
partial_product_5(505) <= '0';
partial_product_5(506) <= '0';
partial_product_5(507) <= '0';
partial_product_5(508) <= '0';
partial_product_5(509) <= '0';
partial_product_5(510) <= '0';
partial_product_5(511) <= '0';
partial_product_5(512) <= '0';
partial_product_6(0) <= '0';
partial_product_6(1) <= '0';
partial_product_6(2) <= '0';
partial_product_6(3) <= '0';
partial_product_6(4) <= '0';
partial_product_6(5) <= '0';
partial_product_6(6) <= '0';
partial_product_6(7) <= '0';
partial_product_6(8) <= '0';
partial_product_6(9) <= '0';
partial_product_6(10) <= '0';
partial_product_6(11) <= '0';
partial_product_6(12) <= '0';
partial_product_6(13) <= '0';
partial_product_6(14) <= '0';
partial_product_6(15) <= '0';
partial_product_6(16) <= '0';
partial_product_6(17) <= '0';
partial_product_6(18) <= '0';
partial_product_6(19) <= '0';
partial_product_6(20) <= '0';
partial_product_6(21) <= '0';
partial_product_6(22) <= '0';
partial_product_6(23) <= '0';
partial_product_6(24) <= '0';
partial_product_6(25) <= '0';
partial_product_6(26) <= '0';
partial_product_6(27) <= '0';
partial_product_6(28) <= '0';
partial_product_6(29) <= '0';
partial_product_6(30) <= '0';
partial_product_6(31) <= '0';
partial_product_6(32) <= '0';
partial_product_6(33) <= '0';
partial_product_6(34) <= '0';
partial_product_6(35) <= '0';
partial_product_6(36) <= '0';
partial_product_6(37) <= '0';
partial_product_6(38) <= '0';
partial_product_6(39) <= '0';
partial_product_6(40) <= '0';
partial_product_6(41) <= '0';
partial_product_6(42) <= '0';
partial_product_6(43) <= '0';
partial_product_6(44) <= '0';
partial_product_6(45) <= '0';
partial_product_6(46) <= '0';
partial_product_6(47) <= '0';
partial_product_6(48) <= '0';
partial_product_6(49) <= '0';
partial_product_6(50) <= '0';
partial_product_6(51) <= '0';
partial_product_6(52) <= '0';
partial_product_6(53) <= '0';
partial_product_6(54) <= '0';
partial_product_6(55) <= '0';
partial_product_6(56) <= '0';
partial_product_6(57) <= '0';
partial_product_6(58) <= '0';
partial_product_6(59) <= '0';
partial_product_6(60) <= '0';
partial_product_6(61) <= '0';
partial_product_6(62) <= '0';
partial_product_6(63) <= '0';
partial_product_6(64) <= '0';
partial_product_6(65) <= '0';
partial_product_6(66) <= '0';
partial_product_6(67) <= '0';
partial_product_6(68) <= temp_mult_20(68);
partial_product_6(69) <= temp_mult_20(69);
partial_product_6(70) <= temp_mult_20(70);
partial_product_6(71) <= temp_mult_20(71);
partial_product_6(72) <= temp_mult_20(72);
partial_product_6(73) <= temp_mult_20(73);
partial_product_6(74) <= temp_mult_20(74);
partial_product_6(75) <= temp_mult_20(75);
partial_product_6(76) <= temp_mult_20(76);
partial_product_6(77) <= temp_mult_20(77);
partial_product_6(78) <= temp_mult_20(78);
partial_product_6(79) <= temp_mult_20(79);
partial_product_6(80) <= temp_mult_20(80);
partial_product_6(81) <= temp_mult_20(81);
partial_product_6(82) <= temp_mult_20(82);
partial_product_6(83) <= temp_mult_20(83);
partial_product_6(84) <= temp_mult_20(84);
partial_product_6(85) <= temp_mult_20(85);
partial_product_6(86) <= temp_mult_20(86);
partial_product_6(87) <= temp_mult_20(87);
partial_product_6(88) <= temp_mult_20(88);
partial_product_6(89) <= temp_mult_20(89);
partial_product_6(90) <= temp_mult_20(90);
partial_product_6(91) <= temp_mult_20(91);
partial_product_6(92) <= temp_mult_20(92);
partial_product_6(93) <= temp_mult_20(93);
partial_product_6(94) <= temp_mult_20(94);
partial_product_6(95) <= temp_mult_20(95);
partial_product_6(96) <= temp_mult_20(96);
partial_product_6(97) <= temp_mult_20(97);
partial_product_6(98) <= temp_mult_20(98);
partial_product_6(99) <= temp_mult_20(99);
partial_product_6(100) <= temp_mult_20(100);
partial_product_6(101) <= temp_mult_20(101);
partial_product_6(102) <= temp_mult_20(102);
partial_product_6(103) <= temp_mult_20(103);
partial_product_6(104) <= temp_mult_20(104);
partial_product_6(105) <= temp_mult_20(105);
partial_product_6(106) <= temp_mult_20(106);
partial_product_6(107) <= temp_mult_20(107);
partial_product_6(108) <= temp_mult_20(108);
partial_product_6(109) <= temp_mult_26(109);
partial_product_6(110) <= temp_mult_26(110);
partial_product_6(111) <= temp_mult_26(111);
partial_product_6(112) <= temp_mult_26(112);
partial_product_6(113) <= temp_mult_26(113);
partial_product_6(114) <= temp_mult_26(114);
partial_product_6(115) <= temp_mult_26(115);
partial_product_6(116) <= temp_mult_26(116);
partial_product_6(117) <= temp_mult_26(117);
partial_product_6(118) <= temp_mult_26(118);
partial_product_6(119) <= temp_mult_26(119);
partial_product_6(120) <= temp_mult_26(120);
partial_product_6(121) <= temp_mult_26(121);
partial_product_6(122) <= temp_mult_26(122);
partial_product_6(123) <= temp_mult_26(123);
partial_product_6(124) <= temp_mult_26(124);
partial_product_6(125) <= temp_mult_26(125);
partial_product_6(126) <= temp_mult_26(126);
partial_product_6(127) <= temp_mult_26(127);
partial_product_6(128) <= temp_mult_26(128);
partial_product_6(129) <= temp_mult_26(129);
partial_product_6(130) <= temp_mult_26(130);
partial_product_6(131) <= temp_mult_26(131);
partial_product_6(132) <= temp_mult_26(132);
partial_product_6(133) <= temp_mult_26(133);
partial_product_6(134) <= temp_mult_26(134);
partial_product_6(135) <= temp_mult_26(135);
partial_product_6(136) <= temp_mult_26(136);
partial_product_6(137) <= temp_mult_26(137);
partial_product_6(138) <= temp_mult_26(138);
partial_product_6(139) <= temp_mult_26(139);
partial_product_6(140) <= temp_mult_26(140);
partial_product_6(141) <= temp_mult_26(141);
partial_product_6(142) <= temp_mult_26(142);
partial_product_6(143) <= temp_mult_26(143);
partial_product_6(144) <= temp_mult_26(144);
partial_product_6(145) <= temp_mult_26(145);
partial_product_6(146) <= temp_mult_26(146);
partial_product_6(147) <= temp_mult_26(147);
partial_product_6(148) <= temp_mult_26(148);
partial_product_6(149) <= temp_mult_26(149);
partial_product_6(150) <= temp_mult_32(150);
partial_product_6(151) <= temp_mult_32(151);
partial_product_6(152) <= temp_mult_32(152);
partial_product_6(153) <= temp_mult_32(153);
partial_product_6(154) <= temp_mult_32(154);
partial_product_6(155) <= temp_mult_32(155);
partial_product_6(156) <= temp_mult_32(156);
partial_product_6(157) <= temp_mult_32(157);
partial_product_6(158) <= temp_mult_32(158);
partial_product_6(159) <= temp_mult_32(159);
partial_product_6(160) <= temp_mult_32(160);
partial_product_6(161) <= temp_mult_32(161);
partial_product_6(162) <= temp_mult_32(162);
partial_product_6(163) <= temp_mult_32(163);
partial_product_6(164) <= temp_mult_32(164);
partial_product_6(165) <= temp_mult_32(165);
partial_product_6(166) <= temp_mult_32(166);
partial_product_6(167) <= temp_mult_32(167);
partial_product_6(168) <= temp_mult_32(168);
partial_product_6(169) <= temp_mult_32(169);
partial_product_6(170) <= temp_mult_32(170);
partial_product_6(171) <= temp_mult_32(171);
partial_product_6(172) <= temp_mult_32(172);
partial_product_6(173) <= temp_mult_32(173);
partial_product_6(174) <= temp_mult_32(174);
partial_product_6(175) <= temp_mult_32(175);
partial_product_6(176) <= temp_mult_32(176);
partial_product_6(177) <= temp_mult_32(177);
partial_product_6(178) <= temp_mult_32(178);
partial_product_6(179) <= temp_mult_32(179);
partial_product_6(180) <= temp_mult_32(180);
partial_product_6(181) <= temp_mult_32(181);
partial_product_6(182) <= temp_mult_32(182);
partial_product_6(183) <= temp_mult_32(183);
partial_product_6(184) <= temp_mult_32(184);
partial_product_6(185) <= temp_mult_32(185);
partial_product_6(186) <= temp_mult_32(186);
partial_product_6(187) <= temp_mult_32(187);
partial_product_6(188) <= temp_mult_32(188);
partial_product_6(189) <= temp_mult_32(189);
partial_product_6(190) <= temp_mult_32(190);
partial_product_6(191) <= temp_mult_38(191);
partial_product_6(192) <= temp_mult_38(192);
partial_product_6(193) <= temp_mult_38(193);
partial_product_6(194) <= temp_mult_38(194);
partial_product_6(195) <= temp_mult_38(195);
partial_product_6(196) <= temp_mult_38(196);
partial_product_6(197) <= temp_mult_38(197);
partial_product_6(198) <= temp_mult_38(198);
partial_product_6(199) <= temp_mult_38(199);
partial_product_6(200) <= temp_mult_38(200);
partial_product_6(201) <= temp_mult_38(201);
partial_product_6(202) <= temp_mult_38(202);
partial_product_6(203) <= temp_mult_38(203);
partial_product_6(204) <= temp_mult_38(204);
partial_product_6(205) <= temp_mult_38(205);
partial_product_6(206) <= temp_mult_38(206);
partial_product_6(207) <= temp_mult_38(207);
partial_product_6(208) <= temp_mult_38(208);
partial_product_6(209) <= temp_mult_38(209);
partial_product_6(210) <= temp_mult_38(210);
partial_product_6(211) <= temp_mult_38(211);
partial_product_6(212) <= temp_mult_38(212);
partial_product_6(213) <= temp_mult_38(213);
partial_product_6(214) <= temp_mult_38(214);
partial_product_6(215) <= temp_mult_38(215);
partial_product_6(216) <= temp_mult_38(216);
partial_product_6(217) <= temp_mult_38(217);
partial_product_6(218) <= temp_mult_38(218);
partial_product_6(219) <= temp_mult_38(219);
partial_product_6(220) <= temp_mult_38(220);
partial_product_6(221) <= temp_mult_38(221);
partial_product_6(222) <= temp_mult_38(222);
partial_product_6(223) <= temp_mult_38(223);
partial_product_6(224) <= temp_mult_38(224);
partial_product_6(225) <= temp_mult_38(225);
partial_product_6(226) <= temp_mult_38(226);
partial_product_6(227) <= temp_mult_38(227);
partial_product_6(228) <= temp_mult_38(228);
partial_product_6(229) <= temp_mult_38(229);
partial_product_6(230) <= temp_mult_38(230);
partial_product_6(231) <= temp_mult_38(231);
partial_product_6(232) <= temp_mult_112(232);
partial_product_6(233) <= temp_mult_112(233);
partial_product_6(234) <= temp_mult_112(234);
partial_product_6(235) <= temp_mult_112(235);
partial_product_6(236) <= temp_mult_112(236);
partial_product_6(237) <= temp_mult_112(237);
partial_product_6(238) <= temp_mult_112(238);
partial_product_6(239) <= temp_mult_112(239);
partial_product_6(240) <= temp_mult_112(240);
partial_product_6(241) <= temp_mult_112(241);
partial_product_6(242) <= temp_mult_112(242);
partial_product_6(243) <= temp_mult_112(243);
partial_product_6(244) <= temp_mult_112(244);
partial_product_6(245) <= temp_mult_112(245);
partial_product_6(246) <= temp_mult_112(246);
partial_product_6(247) <= temp_mult_112(247);
partial_product_6(248) <= temp_mult_112(248);
partial_product_6(249) <= temp_mult_112(249);
partial_product_6(250) <= temp_mult_112(250);
partial_product_6(251) <= temp_mult_112(251);
partial_product_6(252) <= temp_mult_112(252);
partial_product_6(253) <= temp_mult_112(253);
partial_product_6(254) <= temp_mult_112(254);
partial_product_6(255) <= temp_mult_112(255);
partial_product_6(256) <= temp_mult_112(256);
partial_product_6(257) <= temp_mult_112(257);
partial_product_6(258) <= temp_mult_112(258);
partial_product_6(259) <= temp_mult_112(259);
partial_product_6(260) <= temp_mult_112(260);
partial_product_6(261) <= temp_mult_112(261);
partial_product_6(262) <= temp_mult_112(262);
partial_product_6(263) <= temp_mult_112(263);
partial_product_6(264) <= temp_mult_112(264);
partial_product_6(265) <= temp_mult_112(265);
partial_product_6(266) <= temp_mult_112(266);
partial_product_6(267) <= temp_mult_112(267);
partial_product_6(268) <= temp_mult_112(268);
partial_product_6(269) <= temp_mult_112(269);
partial_product_6(270) <= temp_mult_112(270);
partial_product_6(271) <= temp_mult_112(271);
partial_product_6(272) <= temp_mult_112(272);
partial_product_6(273) <= temp_mult_125(273);
partial_product_6(274) <= temp_mult_125(274);
partial_product_6(275) <= temp_mult_125(275);
partial_product_6(276) <= temp_mult_125(276);
partial_product_6(277) <= temp_mult_125(277);
partial_product_6(278) <= temp_mult_125(278);
partial_product_6(279) <= temp_mult_125(279);
partial_product_6(280) <= temp_mult_125(280);
partial_product_6(281) <= temp_mult_125(281);
partial_product_6(282) <= temp_mult_125(282);
partial_product_6(283) <= temp_mult_125(283);
partial_product_6(284) <= temp_mult_125(284);
partial_product_6(285) <= temp_mult_125(285);
partial_product_6(286) <= temp_mult_125(286);
partial_product_6(287) <= temp_mult_125(287);
partial_product_6(288) <= temp_mult_125(288);
partial_product_6(289) <= temp_mult_125(289);
partial_product_6(290) <= temp_mult_125(290);
partial_product_6(291) <= temp_mult_125(291);
partial_product_6(292) <= temp_mult_125(292);
partial_product_6(293) <= temp_mult_125(293);
partial_product_6(294) <= temp_mult_125(294);
partial_product_6(295) <= temp_mult_125(295);
partial_product_6(296) <= temp_mult_125(296);
partial_product_6(297) <= temp_mult_125(297);
partial_product_6(298) <= temp_mult_125(298);
partial_product_6(299) <= temp_mult_125(299);
partial_product_6(300) <= temp_mult_125(300);
partial_product_6(301) <= temp_mult_125(301);
partial_product_6(302) <= temp_mult_125(302);
partial_product_6(303) <= temp_mult_125(303);
partial_product_6(304) <= temp_mult_125(304);
partial_product_6(305) <= temp_mult_125(305);
partial_product_6(306) <= temp_mult_125(306);
partial_product_6(307) <= temp_mult_125(307);
partial_product_6(308) <= temp_mult_125(308);
partial_product_6(309) <= temp_mult_125(309);
partial_product_6(310) <= temp_mult_125(310);
partial_product_6(311) <= temp_mult_125(311);
partial_product_6(312) <= temp_mult_125(312);
partial_product_6(313) <= temp_mult_125(313);
partial_product_6(314) <= temp_mult_131(314);
partial_product_6(315) <= temp_mult_131(315);
partial_product_6(316) <= temp_mult_131(316);
partial_product_6(317) <= temp_mult_131(317);
partial_product_6(318) <= temp_mult_131(318);
partial_product_6(319) <= temp_mult_131(319);
partial_product_6(320) <= temp_mult_131(320);
partial_product_6(321) <= temp_mult_131(321);
partial_product_6(322) <= temp_mult_131(322);
partial_product_6(323) <= temp_mult_131(323);
partial_product_6(324) <= temp_mult_131(324);
partial_product_6(325) <= temp_mult_131(325);
partial_product_6(326) <= temp_mult_131(326);
partial_product_6(327) <= temp_mult_131(327);
partial_product_6(328) <= temp_mult_131(328);
partial_product_6(329) <= temp_mult_131(329);
partial_product_6(330) <= temp_mult_131(330);
partial_product_6(331) <= temp_mult_131(331);
partial_product_6(332) <= temp_mult_131(332);
partial_product_6(333) <= temp_mult_131(333);
partial_product_6(334) <= temp_mult_131(334);
partial_product_6(335) <= temp_mult_131(335);
partial_product_6(336) <= temp_mult_131(336);
partial_product_6(337) <= temp_mult_131(337);
partial_product_6(338) <= temp_mult_131(338);
partial_product_6(339) <= temp_mult_131(339);
partial_product_6(340) <= temp_mult_131(340);
partial_product_6(341) <= temp_mult_131(341);
partial_product_6(342) <= temp_mult_131(342);
partial_product_6(343) <= temp_mult_131(343);
partial_product_6(344) <= temp_mult_131(344);
partial_product_6(345) <= temp_mult_131(345);
partial_product_6(346) <= temp_mult_131(346);
partial_product_6(347) <= temp_mult_131(347);
partial_product_6(348) <= temp_mult_131(348);
partial_product_6(349) <= temp_mult_131(349);
partial_product_6(350) <= temp_mult_131(350);
partial_product_6(351) <= temp_mult_131(351);
partial_product_6(352) <= temp_mult_131(352);
partial_product_6(353) <= temp_mult_131(353);
partial_product_6(354) <= temp_mult_131(354);
partial_product_6(355) <= temp_mult_137(355);
partial_product_6(356) <= temp_mult_137(356);
partial_product_6(357) <= temp_mult_137(357);
partial_product_6(358) <= temp_mult_137(358);
partial_product_6(359) <= temp_mult_137(359);
partial_product_6(360) <= temp_mult_137(360);
partial_product_6(361) <= temp_mult_137(361);
partial_product_6(362) <= temp_mult_137(362);
partial_product_6(363) <= temp_mult_137(363);
partial_product_6(364) <= temp_mult_137(364);
partial_product_6(365) <= temp_mult_137(365);
partial_product_6(366) <= temp_mult_137(366);
partial_product_6(367) <= temp_mult_137(367);
partial_product_6(368) <= temp_mult_137(368);
partial_product_6(369) <= temp_mult_137(369);
partial_product_6(370) <= temp_mult_137(370);
partial_product_6(371) <= temp_mult_137(371);
partial_product_6(372) <= temp_mult_137(372);
partial_product_6(373) <= temp_mult_137(373);
partial_product_6(374) <= temp_mult_137(374);
partial_product_6(375) <= temp_mult_137(375);
partial_product_6(376) <= temp_mult_137(376);
partial_product_6(377) <= temp_mult_137(377);
partial_product_6(378) <= temp_mult_137(378);
partial_product_6(379) <= temp_mult_137(379);
partial_product_6(380) <= temp_mult_137(380);
partial_product_6(381) <= temp_mult_137(381);
partial_product_6(382) <= temp_mult_137(382);
partial_product_6(383) <= temp_mult_137(383);
partial_product_6(384) <= temp_mult_137(384);
partial_product_6(385) <= temp_mult_137(385);
partial_product_6(386) <= temp_mult_137(386);
partial_product_6(387) <= temp_mult_137(387);
partial_product_6(388) <= temp_mult_137(388);
partial_product_6(389) <= temp_mult_137(389);
partial_product_6(390) <= temp_mult_137(390);
partial_product_6(391) <= temp_mult_137(391);
partial_product_6(392) <= temp_mult_137(392);
partial_product_6(393) <= temp_mult_137(393);
partial_product_6(394) <= temp_mult_137(394);
partial_product_6(395) <= temp_mult_137(395);
partial_product_6(396) <= '0';
partial_product_6(397) <= '0';
partial_product_6(398) <= '0';
partial_product_6(399) <= temp_mult_156(399);
partial_product_6(400) <= temp_mult_156(400);
partial_product_6(401) <= temp_mult_156(401);
partial_product_6(402) <= temp_mult_156(402);
partial_product_6(403) <= temp_mult_156(403);
partial_product_6(404) <= temp_mult_156(404);
partial_product_6(405) <= temp_mult_156(405);
partial_product_6(406) <= temp_mult_156(406);
partial_product_6(407) <= temp_mult_156(407);
partial_product_6(408) <= temp_mult_156(408);
partial_product_6(409) <= temp_mult_156(409);
partial_product_6(410) <= temp_mult_156(410);
partial_product_6(411) <= temp_mult_156(411);
partial_product_6(412) <= temp_mult_156(412);
partial_product_6(413) <= temp_mult_156(413);
partial_product_6(414) <= temp_mult_156(414);
partial_product_6(415) <= temp_mult_156(415);
partial_product_6(416) <= temp_mult_156(416);
partial_product_6(417) <= temp_mult_156(417);
partial_product_6(418) <= temp_mult_156(418);
partial_product_6(419) <= temp_mult_156(419);
partial_product_6(420) <= temp_mult_156(420);
partial_product_6(421) <= temp_mult_156(421);
partial_product_6(422) <= temp_mult_156(422);
partial_product_6(423) <= temp_mult_156(423);
partial_product_6(424) <= temp_mult_156(424);
partial_product_6(425) <= temp_mult_156(425);
partial_product_6(426) <= temp_mult_156(426);
partial_product_6(427) <= temp_mult_156(427);
partial_product_6(428) <= temp_mult_156(428);
partial_product_6(429) <= temp_mult_156(429);
partial_product_6(430) <= temp_mult_156(430);
partial_product_6(431) <= temp_mult_156(431);
partial_product_6(432) <= temp_mult_156(432);
partial_product_6(433) <= temp_mult_156(433);
partial_product_6(434) <= temp_mult_156(434);
partial_product_6(435) <= temp_mult_156(435);
partial_product_6(436) <= temp_mult_156(436);
partial_product_6(437) <= temp_mult_156(437);
partial_product_6(438) <= temp_mult_156(438);
partial_product_6(439) <= temp_mult_156(439);
partial_product_6(440) <= '0';
partial_product_6(441) <= '0';
partial_product_6(442) <= '0';
partial_product_6(443) <= '0';
partial_product_6(444) <= '0';
partial_product_6(445) <= '0';
partial_product_6(446) <= '0';
partial_product_6(447) <= '0';
partial_product_6(448) <= '0';
partial_product_6(449) <= '0';
partial_product_6(450) <= '0';
partial_product_6(451) <= '0';
partial_product_6(452) <= '0';
partial_product_6(453) <= '0';
partial_product_6(454) <= '0';
partial_product_6(455) <= '0';
partial_product_6(456) <= '0';
partial_product_6(457) <= '0';
partial_product_6(458) <= '0';
partial_product_6(459) <= '0';
partial_product_6(460) <= '0';
partial_product_6(461) <= '0';
partial_product_6(462) <= '0';
partial_product_6(463) <= '0';
partial_product_6(464) <= '0';
partial_product_6(465) <= '0';
partial_product_6(466) <= '0';
partial_product_6(467) <= '0';
partial_product_6(468) <= '0';
partial_product_6(469) <= '0';
partial_product_6(470) <= '0';
partial_product_6(471) <= '0';
partial_product_6(472) <= '0';
partial_product_6(473) <= '0';
partial_product_6(474) <= '0';
partial_product_6(475) <= '0';
partial_product_6(476) <= '0';
partial_product_6(477) <= '0';
partial_product_6(478) <= '0';
partial_product_6(479) <= '0';
partial_product_6(480) <= '0';
partial_product_6(481) <= '0';
partial_product_6(482) <= '0';
partial_product_6(483) <= '0';
partial_product_6(484) <= '0';
partial_product_6(485) <= '0';
partial_product_6(486) <= '0';
partial_product_6(487) <= '0';
partial_product_6(488) <= '0';
partial_product_6(489) <= '0';
partial_product_6(490) <= '0';
partial_product_6(491) <= '0';
partial_product_6(492) <= '0';
partial_product_6(493) <= '0';
partial_product_6(494) <= '0';
partial_product_6(495) <= '0';
partial_product_6(496) <= '0';
partial_product_6(497) <= '0';
partial_product_6(498) <= '0';
partial_product_6(499) <= '0';
partial_product_6(500) <= '0';
partial_product_6(501) <= '0';
partial_product_6(502) <= '0';
partial_product_6(503) <= '0';
partial_product_6(504) <= '0';
partial_product_6(505) <= '0';
partial_product_6(506) <= '0';
partial_product_6(507) <= '0';
partial_product_6(508) <= '0';
partial_product_6(509) <= '0';
partial_product_6(510) <= '0';
partial_product_6(511) <= '0';
partial_product_6(512) <= '0';
partial_product_7(0) <= '0';
partial_product_7(1) <= '0';
partial_product_7(2) <= '0';
partial_product_7(3) <= '0';
partial_product_7(4) <= '0';
partial_product_7(5) <= '0';
partial_product_7(6) <= '0';
partial_product_7(7) <= '0';
partial_product_7(8) <= '0';
partial_product_7(9) <= '0';
partial_product_7(10) <= '0';
partial_product_7(11) <= '0';
partial_product_7(12) <= '0';
partial_product_7(13) <= '0';
partial_product_7(14) <= '0';
partial_product_7(15) <= '0';
partial_product_7(16) <= '0';
partial_product_7(17) <= '0';
partial_product_7(18) <= '0';
partial_product_7(19) <= '0';
partial_product_7(20) <= '0';
partial_product_7(21) <= '0';
partial_product_7(22) <= '0';
partial_product_7(23) <= '0';
partial_product_7(24) <= '0';
partial_product_7(25) <= '0';
partial_product_7(26) <= '0';
partial_product_7(27) <= '0';
partial_product_7(28) <= '0';
partial_product_7(29) <= '0';
partial_product_7(30) <= '0';
partial_product_7(31) <= '0';
partial_product_7(32) <= '0';
partial_product_7(33) <= '0';
partial_product_7(34) <= '0';
partial_product_7(35) <= '0';
partial_product_7(36) <= '0';
partial_product_7(37) <= '0';
partial_product_7(38) <= '0';
partial_product_7(39) <= '0';
partial_product_7(40) <= '0';
partial_product_7(41) <= '0';
partial_product_7(42) <= '0';
partial_product_7(43) <= '0';
partial_product_7(44) <= '0';
partial_product_7(45) <= '0';
partial_product_7(46) <= '0';
partial_product_7(47) <= '0';
partial_product_7(48) <= '0';
partial_product_7(49) <= '0';
partial_product_7(50) <= '0';
partial_product_7(51) <= '0';
partial_product_7(52) <= '0';
partial_product_7(53) <= '0';
partial_product_7(54) <= '0';
partial_product_7(55) <= '0';
partial_product_7(56) <= '0';
partial_product_7(57) <= '0';
partial_product_7(58) <= '0';
partial_product_7(59) <= '0';
partial_product_7(60) <= '0';
partial_product_7(61) <= '0';
partial_product_7(62) <= '0';
partial_product_7(63) <= '0';
partial_product_7(64) <= '0';
partial_product_7(65) <= '0';
partial_product_7(66) <= '0';
partial_product_7(67) <= '0';
partial_product_7(68) <= '0';
partial_product_7(69) <= '0';
partial_product_7(70) <= '0';
partial_product_7(71) <= '0';
partial_product_7(72) <= temp_mult_3(72);
partial_product_7(73) <= temp_mult_3(73);
partial_product_7(74) <= temp_mult_3(74);
partial_product_7(75) <= temp_mult_3(75);
partial_product_7(76) <= temp_mult_3(76);
partial_product_7(77) <= temp_mult_3(77);
partial_product_7(78) <= temp_mult_3(78);
partial_product_7(79) <= temp_mult_3(79);
partial_product_7(80) <= temp_mult_3(80);
partial_product_7(81) <= temp_mult_3(81);
partial_product_7(82) <= temp_mult_3(82);
partial_product_7(83) <= temp_mult_3(83);
partial_product_7(84) <= temp_mult_3(84);
partial_product_7(85) <= temp_mult_3(85);
partial_product_7(86) <= temp_mult_3(86);
partial_product_7(87) <= temp_mult_3(87);
partial_product_7(88) <= temp_mult_3(88);
partial_product_7(89) <= temp_mult_3(89);
partial_product_7(90) <= temp_mult_3(90);
partial_product_7(91) <= temp_mult_3(91);
partial_product_7(92) <= temp_mult_3(92);
partial_product_7(93) <= temp_mult_3(93);
partial_product_7(94) <= temp_mult_3(94);
partial_product_7(95) <= temp_mult_3(95);
partial_product_7(96) <= temp_mult_3(96);
partial_product_7(97) <= temp_mult_3(97);
partial_product_7(98) <= temp_mult_3(98);
partial_product_7(99) <= temp_mult_3(99);
partial_product_7(100) <= temp_mult_3(100);
partial_product_7(101) <= temp_mult_3(101);
partial_product_7(102) <= temp_mult_3(102);
partial_product_7(103) <= temp_mult_3(103);
partial_product_7(104) <= temp_mult_3(104);
partial_product_7(105) <= temp_mult_3(105);
partial_product_7(106) <= temp_mult_3(106);
partial_product_7(107) <= temp_mult_3(107);
partial_product_7(108) <= temp_mult_3(108);
partial_product_7(109) <= temp_mult_3(109);
partial_product_7(110) <= temp_mult_3(110);
partial_product_7(111) <= temp_mult_3(111);
partial_product_7(112) <= temp_mult_3(112);
partial_product_7(113) <= temp_mult_9(113);
partial_product_7(114) <= temp_mult_9(114);
partial_product_7(115) <= temp_mult_9(115);
partial_product_7(116) <= temp_mult_9(116);
partial_product_7(117) <= temp_mult_9(117);
partial_product_7(118) <= temp_mult_9(118);
partial_product_7(119) <= temp_mult_9(119);
partial_product_7(120) <= temp_mult_9(120);
partial_product_7(121) <= temp_mult_9(121);
partial_product_7(122) <= temp_mult_9(122);
partial_product_7(123) <= temp_mult_9(123);
partial_product_7(124) <= temp_mult_9(124);
partial_product_7(125) <= temp_mult_9(125);
partial_product_7(126) <= temp_mult_9(126);
partial_product_7(127) <= temp_mult_9(127);
partial_product_7(128) <= temp_mult_9(128);
partial_product_7(129) <= temp_mult_9(129);
partial_product_7(130) <= temp_mult_9(130);
partial_product_7(131) <= temp_mult_9(131);
partial_product_7(132) <= temp_mult_9(132);
partial_product_7(133) <= temp_mult_9(133);
partial_product_7(134) <= temp_mult_9(134);
partial_product_7(135) <= temp_mult_9(135);
partial_product_7(136) <= temp_mult_9(136);
partial_product_7(137) <= temp_mult_9(137);
partial_product_7(138) <= temp_mult_9(138);
partial_product_7(139) <= temp_mult_9(139);
partial_product_7(140) <= temp_mult_9(140);
partial_product_7(141) <= temp_mult_9(141);
partial_product_7(142) <= temp_mult_9(142);
partial_product_7(143) <= temp_mult_9(143);
partial_product_7(144) <= temp_mult_9(144);
partial_product_7(145) <= temp_mult_9(145);
partial_product_7(146) <= temp_mult_9(146);
partial_product_7(147) <= temp_mult_9(147);
partial_product_7(148) <= temp_mult_9(148);
partial_product_7(149) <= temp_mult_9(149);
partial_product_7(150) <= temp_mult_9(150);
partial_product_7(151) <= temp_mult_9(151);
partial_product_7(152) <= temp_mult_9(152);
partial_product_7(153) <= temp_mult_9(153);
partial_product_7(154) <= temp_mult_42(154);
partial_product_7(155) <= temp_mult_42(155);
partial_product_7(156) <= temp_mult_42(156);
partial_product_7(157) <= temp_mult_42(157);
partial_product_7(158) <= temp_mult_42(158);
partial_product_7(159) <= temp_mult_42(159);
partial_product_7(160) <= temp_mult_42(160);
partial_product_7(161) <= temp_mult_42(161);
partial_product_7(162) <= temp_mult_42(162);
partial_product_7(163) <= temp_mult_42(163);
partial_product_7(164) <= temp_mult_42(164);
partial_product_7(165) <= temp_mult_42(165);
partial_product_7(166) <= temp_mult_42(166);
partial_product_7(167) <= temp_mult_42(167);
partial_product_7(168) <= temp_mult_42(168);
partial_product_7(169) <= temp_mult_42(169);
partial_product_7(170) <= temp_mult_42(170);
partial_product_7(171) <= temp_mult_42(171);
partial_product_7(172) <= temp_mult_42(172);
partial_product_7(173) <= temp_mult_42(173);
partial_product_7(174) <= temp_mult_42(174);
partial_product_7(175) <= temp_mult_42(175);
partial_product_7(176) <= temp_mult_42(176);
partial_product_7(177) <= temp_mult_42(177);
partial_product_7(178) <= temp_mult_42(178);
partial_product_7(179) <= temp_mult_42(179);
partial_product_7(180) <= temp_mult_42(180);
partial_product_7(181) <= temp_mult_42(181);
partial_product_7(182) <= temp_mult_42(182);
partial_product_7(183) <= temp_mult_42(183);
partial_product_7(184) <= temp_mult_42(184);
partial_product_7(185) <= temp_mult_42(185);
partial_product_7(186) <= temp_mult_42(186);
partial_product_7(187) <= temp_mult_42(187);
partial_product_7(188) <= temp_mult_42(188);
partial_product_7(189) <= temp_mult_42(189);
partial_product_7(190) <= temp_mult_42(190);
partial_product_7(191) <= temp_mult_42(191);
partial_product_7(192) <= temp_mult_42(192);
partial_product_7(193) <= temp_mult_42(193);
partial_product_7(194) <= temp_mult_42(194);
partial_product_7(195) <= temp_mult_51(195);
partial_product_7(196) <= temp_mult_51(196);
partial_product_7(197) <= temp_mult_51(197);
partial_product_7(198) <= temp_mult_51(198);
partial_product_7(199) <= temp_mult_51(199);
partial_product_7(200) <= temp_mult_51(200);
partial_product_7(201) <= temp_mult_51(201);
partial_product_7(202) <= temp_mult_51(202);
partial_product_7(203) <= temp_mult_51(203);
partial_product_7(204) <= temp_mult_51(204);
partial_product_7(205) <= temp_mult_51(205);
partial_product_7(206) <= temp_mult_51(206);
partial_product_7(207) <= temp_mult_51(207);
partial_product_7(208) <= temp_mult_51(208);
partial_product_7(209) <= temp_mult_51(209);
partial_product_7(210) <= temp_mult_51(210);
partial_product_7(211) <= temp_mult_51(211);
partial_product_7(212) <= temp_mult_51(212);
partial_product_7(213) <= temp_mult_51(213);
partial_product_7(214) <= temp_mult_51(214);
partial_product_7(215) <= temp_mult_51(215);
partial_product_7(216) <= temp_mult_51(216);
partial_product_7(217) <= temp_mult_51(217);
partial_product_7(218) <= temp_mult_51(218);
partial_product_7(219) <= temp_mult_51(219);
partial_product_7(220) <= temp_mult_51(220);
partial_product_7(221) <= temp_mult_51(221);
partial_product_7(222) <= temp_mult_51(222);
partial_product_7(223) <= temp_mult_51(223);
partial_product_7(224) <= temp_mult_51(224);
partial_product_7(225) <= temp_mult_51(225);
partial_product_7(226) <= temp_mult_51(226);
partial_product_7(227) <= temp_mult_51(227);
partial_product_7(228) <= temp_mult_51(228);
partial_product_7(229) <= temp_mult_51(229);
partial_product_7(230) <= temp_mult_51(230);
partial_product_7(231) <= temp_mult_51(231);
partial_product_7(232) <= temp_mult_51(232);
partial_product_7(233) <= temp_mult_51(233);
partial_product_7(234) <= temp_mult_51(234);
partial_product_7(235) <= temp_mult_51(235);
partial_product_7(236) <= temp_mult_60(236);
partial_product_7(237) <= temp_mult_60(237);
partial_product_7(238) <= temp_mult_60(238);
partial_product_7(239) <= temp_mult_60(239);
partial_product_7(240) <= temp_mult_60(240);
partial_product_7(241) <= temp_mult_60(241);
partial_product_7(242) <= temp_mult_60(242);
partial_product_7(243) <= temp_mult_60(243);
partial_product_7(244) <= temp_mult_60(244);
partial_product_7(245) <= temp_mult_60(245);
partial_product_7(246) <= temp_mult_60(246);
partial_product_7(247) <= temp_mult_60(247);
partial_product_7(248) <= temp_mult_60(248);
partial_product_7(249) <= temp_mult_60(249);
partial_product_7(250) <= temp_mult_60(250);
partial_product_7(251) <= temp_mult_60(251);
partial_product_7(252) <= temp_mult_60(252);
partial_product_7(253) <= temp_mult_60(253);
partial_product_7(254) <= temp_mult_60(254);
partial_product_7(255) <= temp_mult_60(255);
partial_product_7(256) <= temp_mult_60(256);
partial_product_7(257) <= temp_mult_60(257);
partial_product_7(258) <= temp_mult_60(258);
partial_product_7(259) <= temp_mult_60(259);
partial_product_7(260) <= temp_mult_60(260);
partial_product_7(261) <= temp_mult_60(261);
partial_product_7(262) <= temp_mult_60(262);
partial_product_7(263) <= temp_mult_60(263);
partial_product_7(264) <= temp_mult_60(264);
partial_product_7(265) <= temp_mult_60(265);
partial_product_7(266) <= temp_mult_60(266);
partial_product_7(267) <= temp_mult_60(267);
partial_product_7(268) <= temp_mult_60(268);
partial_product_7(269) <= temp_mult_60(269);
partial_product_7(270) <= temp_mult_60(270);
partial_product_7(271) <= temp_mult_60(271);
partial_product_7(272) <= temp_mult_60(272);
partial_product_7(273) <= temp_mult_60(273);
partial_product_7(274) <= temp_mult_60(274);
partial_product_7(275) <= temp_mult_60(275);
partial_product_7(276) <= temp_mult_60(276);
partial_product_7(277) <= temp_mult_69(277);
partial_product_7(278) <= temp_mult_69(278);
partial_product_7(279) <= temp_mult_69(279);
partial_product_7(280) <= temp_mult_69(280);
partial_product_7(281) <= temp_mult_69(281);
partial_product_7(282) <= temp_mult_69(282);
partial_product_7(283) <= temp_mult_69(283);
partial_product_7(284) <= temp_mult_69(284);
partial_product_7(285) <= temp_mult_69(285);
partial_product_7(286) <= temp_mult_69(286);
partial_product_7(287) <= temp_mult_69(287);
partial_product_7(288) <= temp_mult_69(288);
partial_product_7(289) <= temp_mult_69(289);
partial_product_7(290) <= temp_mult_69(290);
partial_product_7(291) <= temp_mult_69(291);
partial_product_7(292) <= temp_mult_69(292);
partial_product_7(293) <= temp_mult_69(293);
partial_product_7(294) <= temp_mult_69(294);
partial_product_7(295) <= temp_mult_69(295);
partial_product_7(296) <= temp_mult_69(296);
partial_product_7(297) <= temp_mult_69(297);
partial_product_7(298) <= temp_mult_69(298);
partial_product_7(299) <= temp_mult_69(299);
partial_product_7(300) <= temp_mult_69(300);
partial_product_7(301) <= temp_mult_69(301);
partial_product_7(302) <= temp_mult_69(302);
partial_product_7(303) <= temp_mult_69(303);
partial_product_7(304) <= temp_mult_69(304);
partial_product_7(305) <= temp_mult_69(305);
partial_product_7(306) <= temp_mult_69(306);
partial_product_7(307) <= temp_mult_69(307);
partial_product_7(308) <= temp_mult_69(308);
partial_product_7(309) <= temp_mult_69(309);
partial_product_7(310) <= temp_mult_69(310);
partial_product_7(311) <= temp_mult_69(311);
partial_product_7(312) <= temp_mult_69(312);
partial_product_7(313) <= temp_mult_69(313);
partial_product_7(314) <= temp_mult_69(314);
partial_product_7(315) <= temp_mult_69(315);
partial_product_7(316) <= temp_mult_69(316);
partial_product_7(317) <= temp_mult_69(317);
partial_product_7(318) <= temp_mult_78(318);
partial_product_7(319) <= temp_mult_78(319);
partial_product_7(320) <= temp_mult_78(320);
partial_product_7(321) <= temp_mult_78(321);
partial_product_7(322) <= temp_mult_78(322);
partial_product_7(323) <= temp_mult_78(323);
partial_product_7(324) <= temp_mult_78(324);
partial_product_7(325) <= temp_mult_78(325);
partial_product_7(326) <= temp_mult_78(326);
partial_product_7(327) <= temp_mult_78(327);
partial_product_7(328) <= temp_mult_78(328);
partial_product_7(329) <= temp_mult_78(329);
partial_product_7(330) <= temp_mult_78(330);
partial_product_7(331) <= temp_mult_78(331);
partial_product_7(332) <= temp_mult_78(332);
partial_product_7(333) <= temp_mult_78(333);
partial_product_7(334) <= temp_mult_78(334);
partial_product_7(335) <= temp_mult_78(335);
partial_product_7(336) <= temp_mult_78(336);
partial_product_7(337) <= temp_mult_78(337);
partial_product_7(338) <= temp_mult_78(338);
partial_product_7(339) <= temp_mult_78(339);
partial_product_7(340) <= temp_mult_78(340);
partial_product_7(341) <= temp_mult_78(341);
partial_product_7(342) <= temp_mult_78(342);
partial_product_7(343) <= temp_mult_78(343);
partial_product_7(344) <= temp_mult_78(344);
partial_product_7(345) <= temp_mult_78(345);
partial_product_7(346) <= temp_mult_78(346);
partial_product_7(347) <= temp_mult_78(347);
partial_product_7(348) <= temp_mult_78(348);
partial_product_7(349) <= temp_mult_78(349);
partial_product_7(350) <= temp_mult_78(350);
partial_product_7(351) <= temp_mult_78(351);
partial_product_7(352) <= temp_mult_78(352);
partial_product_7(353) <= temp_mult_78(353);
partial_product_7(354) <= temp_mult_78(354);
partial_product_7(355) <= temp_mult_78(355);
partial_product_7(356) <= temp_mult_78(356);
partial_product_7(357) <= temp_mult_78(357);
partial_product_7(358) <= temp_mult_78(358);
partial_product_7(359) <= '0';
partial_product_7(360) <= '0';
partial_product_7(361) <= '0';
partial_product_7(362) <= '0';
partial_product_7(363) <= '0';
partial_product_7(364) <= '0';
partial_product_7(365) <= temp_mult_146(365);
partial_product_7(366) <= temp_mult_146(366);
partial_product_7(367) <= temp_mult_146(367);
partial_product_7(368) <= temp_mult_146(368);
partial_product_7(369) <= temp_mult_146(369);
partial_product_7(370) <= temp_mult_146(370);
partial_product_7(371) <= temp_mult_146(371);
partial_product_7(372) <= temp_mult_146(372);
partial_product_7(373) <= temp_mult_146(373);
partial_product_7(374) <= temp_mult_146(374);
partial_product_7(375) <= temp_mult_146(375);
partial_product_7(376) <= temp_mult_146(376);
partial_product_7(377) <= temp_mult_146(377);
partial_product_7(378) <= temp_mult_146(378);
partial_product_7(379) <= temp_mult_146(379);
partial_product_7(380) <= temp_mult_146(380);
partial_product_7(381) <= temp_mult_146(381);
partial_product_7(382) <= temp_mult_146(382);
partial_product_7(383) <= temp_mult_146(383);
partial_product_7(384) <= temp_mult_146(384);
partial_product_7(385) <= temp_mult_146(385);
partial_product_7(386) <= temp_mult_146(386);
partial_product_7(387) <= temp_mult_146(387);
partial_product_7(388) <= temp_mult_146(388);
partial_product_7(389) <= temp_mult_146(389);
partial_product_7(390) <= temp_mult_146(390);
partial_product_7(391) <= temp_mult_146(391);
partial_product_7(392) <= temp_mult_146(392);
partial_product_7(393) <= temp_mult_146(393);
partial_product_7(394) <= temp_mult_146(394);
partial_product_7(395) <= temp_mult_146(395);
partial_product_7(396) <= temp_mult_146(396);
partial_product_7(397) <= temp_mult_146(397);
partial_product_7(398) <= temp_mult_146(398);
partial_product_7(399) <= temp_mult_146(399);
partial_product_7(400) <= temp_mult_146(400);
partial_product_7(401) <= temp_mult_146(401);
partial_product_7(402) <= temp_mult_146(402);
partial_product_7(403) <= temp_mult_146(403);
partial_product_7(404) <= temp_mult_146(404);
partial_product_7(405) <= temp_mult_146(405);
partial_product_7(406) <= temp_mult_152(406);
partial_product_7(407) <= temp_mult_152(407);
partial_product_7(408) <= temp_mult_152(408);
partial_product_7(409) <= temp_mult_152(409);
partial_product_7(410) <= temp_mult_152(410);
partial_product_7(411) <= temp_mult_152(411);
partial_product_7(412) <= temp_mult_152(412);
partial_product_7(413) <= temp_mult_152(413);
partial_product_7(414) <= temp_mult_152(414);
partial_product_7(415) <= temp_mult_152(415);
partial_product_7(416) <= temp_mult_152(416);
partial_product_7(417) <= temp_mult_152(417);
partial_product_7(418) <= temp_mult_152(418);
partial_product_7(419) <= temp_mult_152(419);
partial_product_7(420) <= temp_mult_152(420);
partial_product_7(421) <= temp_mult_152(421);
partial_product_7(422) <= temp_mult_152(422);
partial_product_7(423) <= temp_mult_152(423);
partial_product_7(424) <= temp_mult_152(424);
partial_product_7(425) <= temp_mult_152(425);
partial_product_7(426) <= temp_mult_152(426);
partial_product_7(427) <= temp_mult_152(427);
partial_product_7(428) <= temp_mult_152(428);
partial_product_7(429) <= temp_mult_152(429);
partial_product_7(430) <= temp_mult_152(430);
partial_product_7(431) <= temp_mult_152(431);
partial_product_7(432) <= temp_mult_152(432);
partial_product_7(433) <= temp_mult_152(433);
partial_product_7(434) <= temp_mult_152(434);
partial_product_7(435) <= temp_mult_152(435);
partial_product_7(436) <= temp_mult_152(436);
partial_product_7(437) <= temp_mult_152(437);
partial_product_7(438) <= temp_mult_152(438);
partial_product_7(439) <= temp_mult_152(439);
partial_product_7(440) <= temp_mult_152(440);
partial_product_7(441) <= temp_mult_152(441);
partial_product_7(442) <= temp_mult_152(442);
partial_product_7(443) <= temp_mult_152(443);
partial_product_7(444) <= temp_mult_152(444);
partial_product_7(445) <= temp_mult_152(445);
partial_product_7(446) <= temp_mult_152(446);
partial_product_7(447) <= '0';
partial_product_7(448) <= '0';
partial_product_7(449) <= '0';
partial_product_7(450) <= '0';
partial_product_7(451) <= '0';
partial_product_7(452) <= '0';
partial_product_7(453) <= '0';
partial_product_7(454) <= '0';
partial_product_7(455) <= '0';
partial_product_7(456) <= '0';
partial_product_7(457) <= '0';
partial_product_7(458) <= '0';
partial_product_7(459) <= '0';
partial_product_7(460) <= '0';
partial_product_7(461) <= '0';
partial_product_7(462) <= '0';
partial_product_7(463) <= '0';
partial_product_7(464) <= '0';
partial_product_7(465) <= '0';
partial_product_7(466) <= '0';
partial_product_7(467) <= '0';
partial_product_7(468) <= '0';
partial_product_7(469) <= '0';
partial_product_7(470) <= '0';
partial_product_7(471) <= '0';
partial_product_7(472) <= '0';
partial_product_7(473) <= '0';
partial_product_7(474) <= '0';
partial_product_7(475) <= '0';
partial_product_7(476) <= '0';
partial_product_7(477) <= '0';
partial_product_7(478) <= '0';
partial_product_7(479) <= '0';
partial_product_7(480) <= '0';
partial_product_7(481) <= '0';
partial_product_7(482) <= '0';
partial_product_7(483) <= '0';
partial_product_7(484) <= '0';
partial_product_7(485) <= '0';
partial_product_7(486) <= '0';
partial_product_7(487) <= '0';
partial_product_7(488) <= '0';
partial_product_7(489) <= '0';
partial_product_7(490) <= '0';
partial_product_7(491) <= '0';
partial_product_7(492) <= '0';
partial_product_7(493) <= '0';
partial_product_7(494) <= '0';
partial_product_7(495) <= '0';
partial_product_7(496) <= '0';
partial_product_7(497) <= '0';
partial_product_7(498) <= '0';
partial_product_7(499) <= '0';
partial_product_7(500) <= '0';
partial_product_7(501) <= '0';
partial_product_7(502) <= '0';
partial_product_7(503) <= '0';
partial_product_7(504) <= '0';
partial_product_7(505) <= '0';
partial_product_7(506) <= '0';
partial_product_7(507) <= '0';
partial_product_7(508) <= '0';
partial_product_7(509) <= '0';
partial_product_7(510) <= '0';
partial_product_7(511) <= '0';
partial_product_7(512) <= '0';
partial_product_8(0) <= '0';
partial_product_8(1) <= '0';
partial_product_8(2) <= '0';
partial_product_8(3) <= '0';
partial_product_8(4) <= '0';
partial_product_8(5) <= '0';
partial_product_8(6) <= '0';
partial_product_8(7) <= '0';
partial_product_8(8) <= '0';
partial_product_8(9) <= '0';
partial_product_8(10) <= '0';
partial_product_8(11) <= '0';
partial_product_8(12) <= '0';
partial_product_8(13) <= '0';
partial_product_8(14) <= '0';
partial_product_8(15) <= '0';
partial_product_8(16) <= '0';
partial_product_8(17) <= '0';
partial_product_8(18) <= '0';
partial_product_8(19) <= '0';
partial_product_8(20) <= '0';
partial_product_8(21) <= '0';
partial_product_8(22) <= '0';
partial_product_8(23) <= '0';
partial_product_8(24) <= '0';
partial_product_8(25) <= '0';
partial_product_8(26) <= '0';
partial_product_8(27) <= '0';
partial_product_8(28) <= '0';
partial_product_8(29) <= '0';
partial_product_8(30) <= '0';
partial_product_8(31) <= '0';
partial_product_8(32) <= '0';
partial_product_8(33) <= '0';
partial_product_8(34) <= '0';
partial_product_8(35) <= '0';
partial_product_8(36) <= '0';
partial_product_8(37) <= '0';
partial_product_8(38) <= '0';
partial_product_8(39) <= '0';
partial_product_8(40) <= '0';
partial_product_8(41) <= '0';
partial_product_8(42) <= '0';
partial_product_8(43) <= '0';
partial_product_8(44) <= '0';
partial_product_8(45) <= '0';
partial_product_8(46) <= '0';
partial_product_8(47) <= '0';
partial_product_8(48) <= '0';
partial_product_8(49) <= '0';
partial_product_8(50) <= '0';
partial_product_8(51) <= '0';
partial_product_8(52) <= '0';
partial_product_8(53) <= '0';
partial_product_8(54) <= '0';
partial_product_8(55) <= '0';
partial_product_8(56) <= '0';
partial_product_8(57) <= '0';
partial_product_8(58) <= '0';
partial_product_8(59) <= '0';
partial_product_8(60) <= '0';
partial_product_8(61) <= '0';
partial_product_8(62) <= '0';
partial_product_8(63) <= '0';
partial_product_8(64) <= '0';
partial_product_8(65) <= '0';
partial_product_8(66) <= '0';
partial_product_8(67) <= '0';
partial_product_8(68) <= '0';
partial_product_8(69) <= '0';
partial_product_8(70) <= '0';
partial_product_8(71) <= '0';
partial_product_8(72) <= '0';
partial_product_8(73) <= '0';
partial_product_8(74) <= '0';
partial_product_8(75) <= '0';
partial_product_8(76) <= '0';
partial_product_8(77) <= '0';
partial_product_8(78) <= '0';
partial_product_8(79) <= '0';
partial_product_8(80) <= '0';
partial_product_8(81) <= '0';
partial_product_8(82) <= '0';
partial_product_8(83) <= '0';
partial_product_8(84) <= '0';
partial_product_8(85) <= temp_mult_25(85);
partial_product_8(86) <= temp_mult_25(86);
partial_product_8(87) <= temp_mult_25(87);
partial_product_8(88) <= temp_mult_25(88);
partial_product_8(89) <= temp_mult_25(89);
partial_product_8(90) <= temp_mult_25(90);
partial_product_8(91) <= temp_mult_25(91);
partial_product_8(92) <= temp_mult_25(92);
partial_product_8(93) <= temp_mult_25(93);
partial_product_8(94) <= temp_mult_25(94);
partial_product_8(95) <= temp_mult_25(95);
partial_product_8(96) <= temp_mult_25(96);
partial_product_8(97) <= temp_mult_25(97);
partial_product_8(98) <= temp_mult_25(98);
partial_product_8(99) <= temp_mult_25(99);
partial_product_8(100) <= temp_mult_25(100);
partial_product_8(101) <= temp_mult_25(101);
partial_product_8(102) <= temp_mult_25(102);
partial_product_8(103) <= temp_mult_25(103);
partial_product_8(104) <= temp_mult_25(104);
partial_product_8(105) <= temp_mult_25(105);
partial_product_8(106) <= temp_mult_25(106);
partial_product_8(107) <= temp_mult_25(107);
partial_product_8(108) <= temp_mult_25(108);
partial_product_8(109) <= temp_mult_25(109);
partial_product_8(110) <= temp_mult_25(110);
partial_product_8(111) <= temp_mult_25(111);
partial_product_8(112) <= temp_mult_25(112);
partial_product_8(113) <= temp_mult_25(113);
partial_product_8(114) <= temp_mult_25(114);
partial_product_8(115) <= temp_mult_25(115);
partial_product_8(116) <= temp_mult_25(116);
partial_product_8(117) <= temp_mult_25(117);
partial_product_8(118) <= temp_mult_25(118);
partial_product_8(119) <= temp_mult_25(119);
partial_product_8(120) <= temp_mult_25(120);
partial_product_8(121) <= temp_mult_25(121);
partial_product_8(122) <= temp_mult_25(122);
partial_product_8(123) <= temp_mult_25(123);
partial_product_8(124) <= temp_mult_25(124);
partial_product_8(125) <= temp_mult_25(125);
partial_product_8(126) <= temp_mult_31(126);
partial_product_8(127) <= temp_mult_31(127);
partial_product_8(128) <= temp_mult_31(128);
partial_product_8(129) <= temp_mult_31(129);
partial_product_8(130) <= temp_mult_31(130);
partial_product_8(131) <= temp_mult_31(131);
partial_product_8(132) <= temp_mult_31(132);
partial_product_8(133) <= temp_mult_31(133);
partial_product_8(134) <= temp_mult_31(134);
partial_product_8(135) <= temp_mult_31(135);
partial_product_8(136) <= temp_mult_31(136);
partial_product_8(137) <= temp_mult_31(137);
partial_product_8(138) <= temp_mult_31(138);
partial_product_8(139) <= temp_mult_31(139);
partial_product_8(140) <= temp_mult_31(140);
partial_product_8(141) <= temp_mult_31(141);
partial_product_8(142) <= temp_mult_31(142);
partial_product_8(143) <= temp_mult_31(143);
partial_product_8(144) <= temp_mult_31(144);
partial_product_8(145) <= temp_mult_31(145);
partial_product_8(146) <= temp_mult_31(146);
partial_product_8(147) <= temp_mult_31(147);
partial_product_8(148) <= temp_mult_31(148);
partial_product_8(149) <= temp_mult_31(149);
partial_product_8(150) <= temp_mult_31(150);
partial_product_8(151) <= temp_mult_31(151);
partial_product_8(152) <= temp_mult_31(152);
partial_product_8(153) <= temp_mult_31(153);
partial_product_8(154) <= temp_mult_31(154);
partial_product_8(155) <= temp_mult_31(155);
partial_product_8(156) <= temp_mult_31(156);
partial_product_8(157) <= temp_mult_31(157);
partial_product_8(158) <= temp_mult_31(158);
partial_product_8(159) <= temp_mult_31(159);
partial_product_8(160) <= temp_mult_31(160);
partial_product_8(161) <= temp_mult_31(161);
partial_product_8(162) <= temp_mult_31(162);
partial_product_8(163) <= temp_mult_31(163);
partial_product_8(164) <= temp_mult_31(164);
partial_product_8(165) <= temp_mult_31(165);
partial_product_8(166) <= temp_mult_31(166);
partial_product_8(167) <= temp_mult_37(167);
partial_product_8(168) <= temp_mult_37(168);
partial_product_8(169) <= temp_mult_37(169);
partial_product_8(170) <= temp_mult_37(170);
partial_product_8(171) <= temp_mult_37(171);
partial_product_8(172) <= temp_mult_37(172);
partial_product_8(173) <= temp_mult_37(173);
partial_product_8(174) <= temp_mult_37(174);
partial_product_8(175) <= temp_mult_37(175);
partial_product_8(176) <= temp_mult_37(176);
partial_product_8(177) <= temp_mult_37(177);
partial_product_8(178) <= temp_mult_37(178);
partial_product_8(179) <= temp_mult_37(179);
partial_product_8(180) <= temp_mult_37(180);
partial_product_8(181) <= temp_mult_37(181);
partial_product_8(182) <= temp_mult_37(182);
partial_product_8(183) <= temp_mult_37(183);
partial_product_8(184) <= temp_mult_37(184);
partial_product_8(185) <= temp_mult_37(185);
partial_product_8(186) <= temp_mult_37(186);
partial_product_8(187) <= temp_mult_37(187);
partial_product_8(188) <= temp_mult_37(188);
partial_product_8(189) <= temp_mult_37(189);
partial_product_8(190) <= temp_mult_37(190);
partial_product_8(191) <= temp_mult_37(191);
partial_product_8(192) <= temp_mult_37(192);
partial_product_8(193) <= temp_mult_37(193);
partial_product_8(194) <= temp_mult_37(194);
partial_product_8(195) <= temp_mult_37(195);
partial_product_8(196) <= temp_mult_37(196);
partial_product_8(197) <= temp_mult_37(197);
partial_product_8(198) <= temp_mult_37(198);
partial_product_8(199) <= temp_mult_37(199);
partial_product_8(200) <= temp_mult_37(200);
partial_product_8(201) <= temp_mult_37(201);
partial_product_8(202) <= temp_mult_37(202);
partial_product_8(203) <= temp_mult_37(203);
partial_product_8(204) <= temp_mult_37(204);
partial_product_8(205) <= temp_mult_37(205);
partial_product_8(206) <= temp_mult_37(206);
partial_product_8(207) <= temp_mult_37(207);
partial_product_8(208) <= temp_mult_104(208);
partial_product_8(209) <= temp_mult_104(209);
partial_product_8(210) <= temp_mult_104(210);
partial_product_8(211) <= temp_mult_104(211);
partial_product_8(212) <= temp_mult_104(212);
partial_product_8(213) <= temp_mult_104(213);
partial_product_8(214) <= temp_mult_104(214);
partial_product_8(215) <= temp_mult_104(215);
partial_product_8(216) <= temp_mult_104(216);
partial_product_8(217) <= temp_mult_104(217);
partial_product_8(218) <= temp_mult_104(218);
partial_product_8(219) <= temp_mult_104(219);
partial_product_8(220) <= temp_mult_104(220);
partial_product_8(221) <= temp_mult_104(221);
partial_product_8(222) <= temp_mult_104(222);
partial_product_8(223) <= temp_mult_104(223);
partial_product_8(224) <= temp_mult_104(224);
partial_product_8(225) <= temp_mult_104(225);
partial_product_8(226) <= temp_mult_104(226);
partial_product_8(227) <= temp_mult_104(227);
partial_product_8(228) <= temp_mult_104(228);
partial_product_8(229) <= temp_mult_104(229);
partial_product_8(230) <= temp_mult_104(230);
partial_product_8(231) <= temp_mult_104(231);
partial_product_8(232) <= temp_mult_104(232);
partial_product_8(233) <= temp_mult_104(233);
partial_product_8(234) <= temp_mult_104(234);
partial_product_8(235) <= temp_mult_104(235);
partial_product_8(236) <= temp_mult_104(236);
partial_product_8(237) <= temp_mult_104(237);
partial_product_8(238) <= temp_mult_104(238);
partial_product_8(239) <= temp_mult_104(239);
partial_product_8(240) <= temp_mult_104(240);
partial_product_8(241) <= temp_mult_104(241);
partial_product_8(242) <= temp_mult_104(242);
partial_product_8(243) <= temp_mult_104(243);
partial_product_8(244) <= temp_mult_104(244);
partial_product_8(245) <= temp_mult_104(245);
partial_product_8(246) <= temp_mult_104(246);
partial_product_8(247) <= temp_mult_104(247);
partial_product_8(248) <= temp_mult_104(248);
partial_product_8(249) <= temp_mult_113(249);
partial_product_8(250) <= temp_mult_113(250);
partial_product_8(251) <= temp_mult_113(251);
partial_product_8(252) <= temp_mult_113(252);
partial_product_8(253) <= temp_mult_113(253);
partial_product_8(254) <= temp_mult_113(254);
partial_product_8(255) <= temp_mult_113(255);
partial_product_8(256) <= temp_mult_113(256);
partial_product_8(257) <= temp_mult_113(257);
partial_product_8(258) <= temp_mult_113(258);
partial_product_8(259) <= temp_mult_113(259);
partial_product_8(260) <= temp_mult_113(260);
partial_product_8(261) <= temp_mult_113(261);
partial_product_8(262) <= temp_mult_113(262);
partial_product_8(263) <= temp_mult_113(263);
partial_product_8(264) <= temp_mult_113(264);
partial_product_8(265) <= temp_mult_113(265);
partial_product_8(266) <= temp_mult_113(266);
partial_product_8(267) <= temp_mult_113(267);
partial_product_8(268) <= temp_mult_113(268);
partial_product_8(269) <= temp_mult_113(269);
partial_product_8(270) <= temp_mult_113(270);
partial_product_8(271) <= temp_mult_113(271);
partial_product_8(272) <= temp_mult_113(272);
partial_product_8(273) <= temp_mult_113(273);
partial_product_8(274) <= temp_mult_113(274);
partial_product_8(275) <= temp_mult_113(275);
partial_product_8(276) <= temp_mult_113(276);
partial_product_8(277) <= temp_mult_113(277);
partial_product_8(278) <= temp_mult_113(278);
partial_product_8(279) <= temp_mult_113(279);
partial_product_8(280) <= temp_mult_113(280);
partial_product_8(281) <= temp_mult_113(281);
partial_product_8(282) <= temp_mult_113(282);
partial_product_8(283) <= temp_mult_113(283);
partial_product_8(284) <= temp_mult_113(284);
partial_product_8(285) <= temp_mult_113(285);
partial_product_8(286) <= temp_mult_113(286);
partial_product_8(287) <= temp_mult_113(287);
partial_product_8(288) <= temp_mult_113(288);
partial_product_8(289) <= temp_mult_113(289);
partial_product_8(290) <= temp_mult_130(290);
partial_product_8(291) <= temp_mult_130(291);
partial_product_8(292) <= temp_mult_130(292);
partial_product_8(293) <= temp_mult_130(293);
partial_product_8(294) <= temp_mult_130(294);
partial_product_8(295) <= temp_mult_130(295);
partial_product_8(296) <= temp_mult_130(296);
partial_product_8(297) <= temp_mult_130(297);
partial_product_8(298) <= temp_mult_130(298);
partial_product_8(299) <= temp_mult_130(299);
partial_product_8(300) <= temp_mult_130(300);
partial_product_8(301) <= temp_mult_130(301);
partial_product_8(302) <= temp_mult_130(302);
partial_product_8(303) <= temp_mult_130(303);
partial_product_8(304) <= temp_mult_130(304);
partial_product_8(305) <= temp_mult_130(305);
partial_product_8(306) <= temp_mult_130(306);
partial_product_8(307) <= temp_mult_130(307);
partial_product_8(308) <= temp_mult_130(308);
partial_product_8(309) <= temp_mult_130(309);
partial_product_8(310) <= temp_mult_130(310);
partial_product_8(311) <= temp_mult_130(311);
partial_product_8(312) <= temp_mult_130(312);
partial_product_8(313) <= temp_mult_130(313);
partial_product_8(314) <= temp_mult_130(314);
partial_product_8(315) <= temp_mult_130(315);
partial_product_8(316) <= temp_mult_130(316);
partial_product_8(317) <= temp_mult_130(317);
partial_product_8(318) <= temp_mult_130(318);
partial_product_8(319) <= temp_mult_130(319);
partial_product_8(320) <= temp_mult_130(320);
partial_product_8(321) <= temp_mult_130(321);
partial_product_8(322) <= temp_mult_130(322);
partial_product_8(323) <= temp_mult_130(323);
partial_product_8(324) <= temp_mult_130(324);
partial_product_8(325) <= temp_mult_130(325);
partial_product_8(326) <= temp_mult_130(326);
partial_product_8(327) <= temp_mult_130(327);
partial_product_8(328) <= temp_mult_130(328);
partial_product_8(329) <= temp_mult_130(329);
partial_product_8(330) <= temp_mult_130(330);
partial_product_8(331) <= temp_mult_136(331);
partial_product_8(332) <= temp_mult_136(332);
partial_product_8(333) <= temp_mult_136(333);
partial_product_8(334) <= temp_mult_136(334);
partial_product_8(335) <= temp_mult_136(335);
partial_product_8(336) <= temp_mult_136(336);
partial_product_8(337) <= temp_mult_136(337);
partial_product_8(338) <= temp_mult_136(338);
partial_product_8(339) <= temp_mult_136(339);
partial_product_8(340) <= temp_mult_136(340);
partial_product_8(341) <= temp_mult_136(341);
partial_product_8(342) <= temp_mult_136(342);
partial_product_8(343) <= temp_mult_136(343);
partial_product_8(344) <= temp_mult_136(344);
partial_product_8(345) <= temp_mult_136(345);
partial_product_8(346) <= temp_mult_136(346);
partial_product_8(347) <= temp_mult_136(347);
partial_product_8(348) <= temp_mult_136(348);
partial_product_8(349) <= temp_mult_136(349);
partial_product_8(350) <= temp_mult_136(350);
partial_product_8(351) <= temp_mult_136(351);
partial_product_8(352) <= temp_mult_136(352);
partial_product_8(353) <= temp_mult_136(353);
partial_product_8(354) <= temp_mult_136(354);
partial_product_8(355) <= temp_mult_136(355);
partial_product_8(356) <= temp_mult_136(356);
partial_product_8(357) <= temp_mult_136(357);
partial_product_8(358) <= temp_mult_136(358);
partial_product_8(359) <= temp_mult_136(359);
partial_product_8(360) <= temp_mult_136(360);
partial_product_8(361) <= temp_mult_136(361);
partial_product_8(362) <= temp_mult_136(362);
partial_product_8(363) <= temp_mult_136(363);
partial_product_8(364) <= temp_mult_136(364);
partial_product_8(365) <= temp_mult_136(365);
partial_product_8(366) <= temp_mult_136(366);
partial_product_8(367) <= temp_mult_136(367);
partial_product_8(368) <= temp_mult_136(368);
partial_product_8(369) <= temp_mult_136(369);
partial_product_8(370) <= temp_mult_136(370);
partial_product_8(371) <= temp_mult_136(371);
partial_product_8(372) <= temp_mult_142(372);
partial_product_8(373) <= temp_mult_142(373);
partial_product_8(374) <= temp_mult_142(374);
partial_product_8(375) <= temp_mult_142(375);
partial_product_8(376) <= temp_mult_142(376);
partial_product_8(377) <= temp_mult_142(377);
partial_product_8(378) <= temp_mult_142(378);
partial_product_8(379) <= temp_mult_142(379);
partial_product_8(380) <= temp_mult_142(380);
partial_product_8(381) <= temp_mult_142(381);
partial_product_8(382) <= temp_mult_142(382);
partial_product_8(383) <= temp_mult_142(383);
partial_product_8(384) <= temp_mult_142(384);
partial_product_8(385) <= temp_mult_142(385);
partial_product_8(386) <= temp_mult_142(386);
partial_product_8(387) <= temp_mult_142(387);
partial_product_8(388) <= temp_mult_142(388);
partial_product_8(389) <= temp_mult_142(389);
partial_product_8(390) <= temp_mult_142(390);
partial_product_8(391) <= temp_mult_142(391);
partial_product_8(392) <= temp_mult_142(392);
partial_product_8(393) <= temp_mult_142(393);
partial_product_8(394) <= temp_mult_142(394);
partial_product_8(395) <= temp_mult_142(395);
partial_product_8(396) <= temp_mult_142(396);
partial_product_8(397) <= temp_mult_142(397);
partial_product_8(398) <= temp_mult_142(398);
partial_product_8(399) <= temp_mult_142(399);
partial_product_8(400) <= temp_mult_142(400);
partial_product_8(401) <= temp_mult_142(401);
partial_product_8(402) <= temp_mult_142(402);
partial_product_8(403) <= temp_mult_142(403);
partial_product_8(404) <= temp_mult_142(404);
partial_product_8(405) <= temp_mult_142(405);
partial_product_8(406) <= temp_mult_142(406);
partial_product_8(407) <= temp_mult_142(407);
partial_product_8(408) <= temp_mult_142(408);
partial_product_8(409) <= temp_mult_142(409);
partial_product_8(410) <= temp_mult_142(410);
partial_product_8(411) <= temp_mult_142(411);
partial_product_8(412) <= temp_mult_142(412);
partial_product_8(413) <= '0';
partial_product_8(414) <= '0';
partial_product_8(415) <= '0';
partial_product_8(416) <= '0';
partial_product_8(417) <= '0';
partial_product_8(418) <= '0';
partial_product_8(419) <= '0';
partial_product_8(420) <= '0';
partial_product_8(421) <= '0';
partial_product_8(422) <= '0';
partial_product_8(423) <= '0';
partial_product_8(424) <= '0';
partial_product_8(425) <= '0';
partial_product_8(426) <= '0';
partial_product_8(427) <= '0';
partial_product_8(428) <= '0';
partial_product_8(429) <= '0';
partial_product_8(430) <= '0';
partial_product_8(431) <= '0';
partial_product_8(432) <= '0';
partial_product_8(433) <= '0';
partial_product_8(434) <= '0';
partial_product_8(435) <= '0';
partial_product_8(436) <= '0';
partial_product_8(437) <= '0';
partial_product_8(438) <= '0';
partial_product_8(439) <= '0';
partial_product_8(440) <= '0';
partial_product_8(441) <= '0';
partial_product_8(442) <= '0';
partial_product_8(443) <= '0';
partial_product_8(444) <= '0';
partial_product_8(445) <= '0';
partial_product_8(446) <= '0';
partial_product_8(447) <= '0';
partial_product_8(448) <= '0';
partial_product_8(449) <= '0';
partial_product_8(450) <= '0';
partial_product_8(451) <= '0';
partial_product_8(452) <= '0';
partial_product_8(453) <= '0';
partial_product_8(454) <= '0';
partial_product_8(455) <= '0';
partial_product_8(456) <= '0';
partial_product_8(457) <= '0';
partial_product_8(458) <= '0';
partial_product_8(459) <= '0';
partial_product_8(460) <= '0';
partial_product_8(461) <= '0';
partial_product_8(462) <= '0';
partial_product_8(463) <= '0';
partial_product_8(464) <= '0';
partial_product_8(465) <= '0';
partial_product_8(466) <= '0';
partial_product_8(467) <= '0';
partial_product_8(468) <= '0';
partial_product_8(469) <= '0';
partial_product_8(470) <= '0';
partial_product_8(471) <= '0';
partial_product_8(472) <= '0';
partial_product_8(473) <= '0';
partial_product_8(474) <= '0';
partial_product_8(475) <= '0';
partial_product_8(476) <= '0';
partial_product_8(477) <= '0';
partial_product_8(478) <= '0';
partial_product_8(479) <= '0';
partial_product_8(480) <= '0';
partial_product_8(481) <= '0';
partial_product_8(482) <= '0';
partial_product_8(483) <= '0';
partial_product_8(484) <= '0';
partial_product_8(485) <= '0';
partial_product_8(486) <= '0';
partial_product_8(487) <= '0';
partial_product_8(488) <= '0';
partial_product_8(489) <= '0';
partial_product_8(490) <= '0';
partial_product_8(491) <= '0';
partial_product_8(492) <= '0';
partial_product_8(493) <= '0';
partial_product_8(494) <= '0';
partial_product_8(495) <= '0';
partial_product_8(496) <= '0';
partial_product_8(497) <= '0';
partial_product_8(498) <= '0';
partial_product_8(499) <= '0';
partial_product_8(500) <= '0';
partial_product_8(501) <= '0';
partial_product_8(502) <= '0';
partial_product_8(503) <= '0';
partial_product_8(504) <= '0';
partial_product_8(505) <= '0';
partial_product_8(506) <= '0';
partial_product_8(507) <= '0';
partial_product_8(508) <= '0';
partial_product_8(509) <= '0';
partial_product_8(510) <= '0';
partial_product_8(511) <= '0';
partial_product_8(512) <= '0';
partial_product_9(0) <= '0';
partial_product_9(1) <= '0';
partial_product_9(2) <= '0';
partial_product_9(3) <= '0';
partial_product_9(4) <= '0';
partial_product_9(5) <= '0';
partial_product_9(6) <= '0';
partial_product_9(7) <= '0';
partial_product_9(8) <= '0';
partial_product_9(9) <= '0';
partial_product_9(10) <= '0';
partial_product_9(11) <= '0';
partial_product_9(12) <= '0';
partial_product_9(13) <= '0';
partial_product_9(14) <= '0';
partial_product_9(15) <= '0';
partial_product_9(16) <= '0';
partial_product_9(17) <= '0';
partial_product_9(18) <= '0';
partial_product_9(19) <= '0';
partial_product_9(20) <= '0';
partial_product_9(21) <= '0';
partial_product_9(22) <= '0';
partial_product_9(23) <= '0';
partial_product_9(24) <= '0';
partial_product_9(25) <= '0';
partial_product_9(26) <= '0';
partial_product_9(27) <= '0';
partial_product_9(28) <= '0';
partial_product_9(29) <= '0';
partial_product_9(30) <= '0';
partial_product_9(31) <= '0';
partial_product_9(32) <= '0';
partial_product_9(33) <= '0';
partial_product_9(34) <= '0';
partial_product_9(35) <= '0';
partial_product_9(36) <= '0';
partial_product_9(37) <= '0';
partial_product_9(38) <= '0';
partial_product_9(39) <= '0';
partial_product_9(40) <= '0';
partial_product_9(41) <= '0';
partial_product_9(42) <= '0';
partial_product_9(43) <= '0';
partial_product_9(44) <= '0';
partial_product_9(45) <= '0';
partial_product_9(46) <= '0';
partial_product_9(47) <= '0';
partial_product_9(48) <= '0';
partial_product_9(49) <= '0';
partial_product_9(50) <= '0';
partial_product_9(51) <= '0';
partial_product_9(52) <= '0';
partial_product_9(53) <= '0';
partial_product_9(54) <= '0';
partial_product_9(55) <= '0';
partial_product_9(56) <= '0';
partial_product_9(57) <= '0';
partial_product_9(58) <= '0';
partial_product_9(59) <= '0';
partial_product_9(60) <= '0';
partial_product_9(61) <= '0';
partial_product_9(62) <= '0';
partial_product_9(63) <= '0';
partial_product_9(64) <= '0';
partial_product_9(65) <= '0';
partial_product_9(66) <= '0';
partial_product_9(67) <= '0';
partial_product_9(68) <= '0';
partial_product_9(69) <= '0';
partial_product_9(70) <= '0';
partial_product_9(71) <= '0';
partial_product_9(72) <= '0';
partial_product_9(73) <= '0';
partial_product_9(74) <= '0';
partial_product_9(75) <= '0';
partial_product_9(76) <= '0';
partial_product_9(77) <= '0';
partial_product_9(78) <= '0';
partial_product_9(79) <= '0';
partial_product_9(80) <= '0';
partial_product_9(81) <= '0';
partial_product_9(82) <= '0';
partial_product_9(83) <= '0';
partial_product_9(84) <= '0';
partial_product_9(85) <= '0';
partial_product_9(86) <= '0';
partial_product_9(87) <= '0';
partial_product_9(88) <= '0';
partial_product_9(89) <= '0';
partial_product_9(90) <= '0';
partial_product_9(91) <= '0';
partial_product_9(92) <= '0';
partial_product_9(93) <= '0';
partial_product_9(94) <= '0';
partial_product_9(95) <= '0';
partial_product_9(96) <= temp_mult_4(96);
partial_product_9(97) <= temp_mult_4(97);
partial_product_9(98) <= temp_mult_4(98);
partial_product_9(99) <= temp_mult_4(99);
partial_product_9(100) <= temp_mult_4(100);
partial_product_9(101) <= temp_mult_4(101);
partial_product_9(102) <= temp_mult_4(102);
partial_product_9(103) <= temp_mult_4(103);
partial_product_9(104) <= temp_mult_4(104);
partial_product_9(105) <= temp_mult_4(105);
partial_product_9(106) <= temp_mult_4(106);
partial_product_9(107) <= temp_mult_4(107);
partial_product_9(108) <= temp_mult_4(108);
partial_product_9(109) <= temp_mult_4(109);
partial_product_9(110) <= temp_mult_4(110);
partial_product_9(111) <= temp_mult_4(111);
partial_product_9(112) <= temp_mult_4(112);
partial_product_9(113) <= temp_mult_4(113);
partial_product_9(114) <= temp_mult_4(114);
partial_product_9(115) <= temp_mult_4(115);
partial_product_9(116) <= temp_mult_4(116);
partial_product_9(117) <= temp_mult_4(117);
partial_product_9(118) <= temp_mult_4(118);
partial_product_9(119) <= temp_mult_4(119);
partial_product_9(120) <= temp_mult_4(120);
partial_product_9(121) <= temp_mult_4(121);
partial_product_9(122) <= temp_mult_4(122);
partial_product_9(123) <= temp_mult_4(123);
partial_product_9(124) <= temp_mult_4(124);
partial_product_9(125) <= temp_mult_4(125);
partial_product_9(126) <= temp_mult_4(126);
partial_product_9(127) <= temp_mult_4(127);
partial_product_9(128) <= temp_mult_4(128);
partial_product_9(129) <= temp_mult_4(129);
partial_product_9(130) <= temp_mult_4(130);
partial_product_9(131) <= temp_mult_4(131);
partial_product_9(132) <= temp_mult_4(132);
partial_product_9(133) <= temp_mult_4(133);
partial_product_9(134) <= temp_mult_4(134);
partial_product_9(135) <= temp_mult_4(135);
partial_product_9(136) <= temp_mult_4(136);
partial_product_9(137) <= temp_mult_41(137);
partial_product_9(138) <= temp_mult_41(138);
partial_product_9(139) <= temp_mult_41(139);
partial_product_9(140) <= temp_mult_41(140);
partial_product_9(141) <= temp_mult_41(141);
partial_product_9(142) <= temp_mult_41(142);
partial_product_9(143) <= temp_mult_41(143);
partial_product_9(144) <= temp_mult_41(144);
partial_product_9(145) <= temp_mult_41(145);
partial_product_9(146) <= temp_mult_41(146);
partial_product_9(147) <= temp_mult_41(147);
partial_product_9(148) <= temp_mult_41(148);
partial_product_9(149) <= temp_mult_41(149);
partial_product_9(150) <= temp_mult_41(150);
partial_product_9(151) <= temp_mult_41(151);
partial_product_9(152) <= temp_mult_41(152);
partial_product_9(153) <= temp_mult_41(153);
partial_product_9(154) <= temp_mult_41(154);
partial_product_9(155) <= temp_mult_41(155);
partial_product_9(156) <= temp_mult_41(156);
partial_product_9(157) <= temp_mult_41(157);
partial_product_9(158) <= temp_mult_41(158);
partial_product_9(159) <= temp_mult_41(159);
partial_product_9(160) <= temp_mult_41(160);
partial_product_9(161) <= temp_mult_41(161);
partial_product_9(162) <= temp_mult_41(162);
partial_product_9(163) <= temp_mult_41(163);
partial_product_9(164) <= temp_mult_41(164);
partial_product_9(165) <= temp_mult_41(165);
partial_product_9(166) <= temp_mult_41(166);
partial_product_9(167) <= temp_mult_41(167);
partial_product_9(168) <= temp_mult_41(168);
partial_product_9(169) <= temp_mult_41(169);
partial_product_9(170) <= temp_mult_41(170);
partial_product_9(171) <= temp_mult_41(171);
partial_product_9(172) <= temp_mult_41(172);
partial_product_9(173) <= temp_mult_41(173);
partial_product_9(174) <= temp_mult_41(174);
partial_product_9(175) <= temp_mult_41(175);
partial_product_9(176) <= temp_mult_41(176);
partial_product_9(177) <= temp_mult_41(177);
partial_product_9(178) <= temp_mult_50(178);
partial_product_9(179) <= temp_mult_50(179);
partial_product_9(180) <= temp_mult_50(180);
partial_product_9(181) <= temp_mult_50(181);
partial_product_9(182) <= temp_mult_50(182);
partial_product_9(183) <= temp_mult_50(183);
partial_product_9(184) <= temp_mult_50(184);
partial_product_9(185) <= temp_mult_50(185);
partial_product_9(186) <= temp_mult_50(186);
partial_product_9(187) <= temp_mult_50(187);
partial_product_9(188) <= temp_mult_50(188);
partial_product_9(189) <= temp_mult_50(189);
partial_product_9(190) <= temp_mult_50(190);
partial_product_9(191) <= temp_mult_50(191);
partial_product_9(192) <= temp_mult_50(192);
partial_product_9(193) <= temp_mult_50(193);
partial_product_9(194) <= temp_mult_50(194);
partial_product_9(195) <= temp_mult_50(195);
partial_product_9(196) <= temp_mult_50(196);
partial_product_9(197) <= temp_mult_50(197);
partial_product_9(198) <= temp_mult_50(198);
partial_product_9(199) <= temp_mult_50(199);
partial_product_9(200) <= temp_mult_50(200);
partial_product_9(201) <= temp_mult_50(201);
partial_product_9(202) <= temp_mult_50(202);
partial_product_9(203) <= temp_mult_50(203);
partial_product_9(204) <= temp_mult_50(204);
partial_product_9(205) <= temp_mult_50(205);
partial_product_9(206) <= temp_mult_50(206);
partial_product_9(207) <= temp_mult_50(207);
partial_product_9(208) <= temp_mult_50(208);
partial_product_9(209) <= temp_mult_50(209);
partial_product_9(210) <= temp_mult_50(210);
partial_product_9(211) <= temp_mult_50(211);
partial_product_9(212) <= temp_mult_50(212);
partial_product_9(213) <= temp_mult_50(213);
partial_product_9(214) <= temp_mult_50(214);
partial_product_9(215) <= temp_mult_50(215);
partial_product_9(216) <= temp_mult_50(216);
partial_product_9(217) <= temp_mult_50(217);
partial_product_9(218) <= temp_mult_50(218);
partial_product_9(219) <= temp_mult_59(219);
partial_product_9(220) <= temp_mult_59(220);
partial_product_9(221) <= temp_mult_59(221);
partial_product_9(222) <= temp_mult_59(222);
partial_product_9(223) <= temp_mult_59(223);
partial_product_9(224) <= temp_mult_59(224);
partial_product_9(225) <= temp_mult_59(225);
partial_product_9(226) <= temp_mult_59(226);
partial_product_9(227) <= temp_mult_59(227);
partial_product_9(228) <= temp_mult_59(228);
partial_product_9(229) <= temp_mult_59(229);
partial_product_9(230) <= temp_mult_59(230);
partial_product_9(231) <= temp_mult_59(231);
partial_product_9(232) <= temp_mult_59(232);
partial_product_9(233) <= temp_mult_59(233);
partial_product_9(234) <= temp_mult_59(234);
partial_product_9(235) <= temp_mult_59(235);
partial_product_9(236) <= temp_mult_59(236);
partial_product_9(237) <= temp_mult_59(237);
partial_product_9(238) <= temp_mult_59(238);
partial_product_9(239) <= temp_mult_59(239);
partial_product_9(240) <= temp_mult_59(240);
partial_product_9(241) <= temp_mult_59(241);
partial_product_9(242) <= temp_mult_59(242);
partial_product_9(243) <= temp_mult_59(243);
partial_product_9(244) <= temp_mult_59(244);
partial_product_9(245) <= temp_mult_59(245);
partial_product_9(246) <= temp_mult_59(246);
partial_product_9(247) <= temp_mult_59(247);
partial_product_9(248) <= temp_mult_59(248);
partial_product_9(249) <= temp_mult_59(249);
partial_product_9(250) <= temp_mult_59(250);
partial_product_9(251) <= temp_mult_59(251);
partial_product_9(252) <= temp_mult_59(252);
partial_product_9(253) <= temp_mult_59(253);
partial_product_9(254) <= temp_mult_59(254);
partial_product_9(255) <= temp_mult_59(255);
partial_product_9(256) <= temp_mult_59(256);
partial_product_9(257) <= temp_mult_59(257);
partial_product_9(258) <= temp_mult_59(258);
partial_product_9(259) <= temp_mult_59(259);
partial_product_9(260) <= temp_mult_68(260);
partial_product_9(261) <= temp_mult_68(261);
partial_product_9(262) <= temp_mult_68(262);
partial_product_9(263) <= temp_mult_68(263);
partial_product_9(264) <= temp_mult_68(264);
partial_product_9(265) <= temp_mult_68(265);
partial_product_9(266) <= temp_mult_68(266);
partial_product_9(267) <= temp_mult_68(267);
partial_product_9(268) <= temp_mult_68(268);
partial_product_9(269) <= temp_mult_68(269);
partial_product_9(270) <= temp_mult_68(270);
partial_product_9(271) <= temp_mult_68(271);
partial_product_9(272) <= temp_mult_68(272);
partial_product_9(273) <= temp_mult_68(273);
partial_product_9(274) <= temp_mult_68(274);
partial_product_9(275) <= temp_mult_68(275);
partial_product_9(276) <= temp_mult_68(276);
partial_product_9(277) <= temp_mult_68(277);
partial_product_9(278) <= temp_mult_68(278);
partial_product_9(279) <= temp_mult_68(279);
partial_product_9(280) <= temp_mult_68(280);
partial_product_9(281) <= temp_mult_68(281);
partial_product_9(282) <= temp_mult_68(282);
partial_product_9(283) <= temp_mult_68(283);
partial_product_9(284) <= temp_mult_68(284);
partial_product_9(285) <= temp_mult_68(285);
partial_product_9(286) <= temp_mult_68(286);
partial_product_9(287) <= temp_mult_68(287);
partial_product_9(288) <= temp_mult_68(288);
partial_product_9(289) <= temp_mult_68(289);
partial_product_9(290) <= temp_mult_68(290);
partial_product_9(291) <= temp_mult_68(291);
partial_product_9(292) <= temp_mult_68(292);
partial_product_9(293) <= temp_mult_68(293);
partial_product_9(294) <= temp_mult_68(294);
partial_product_9(295) <= temp_mult_68(295);
partial_product_9(296) <= temp_mult_68(296);
partial_product_9(297) <= temp_mult_68(297);
partial_product_9(298) <= temp_mult_68(298);
partial_product_9(299) <= temp_mult_68(299);
partial_product_9(300) <= temp_mult_68(300);
partial_product_9(301) <= temp_mult_77(301);
partial_product_9(302) <= temp_mult_77(302);
partial_product_9(303) <= temp_mult_77(303);
partial_product_9(304) <= temp_mult_77(304);
partial_product_9(305) <= temp_mult_77(305);
partial_product_9(306) <= temp_mult_77(306);
partial_product_9(307) <= temp_mult_77(307);
partial_product_9(308) <= temp_mult_77(308);
partial_product_9(309) <= temp_mult_77(309);
partial_product_9(310) <= temp_mult_77(310);
partial_product_9(311) <= temp_mult_77(311);
partial_product_9(312) <= temp_mult_77(312);
partial_product_9(313) <= temp_mult_77(313);
partial_product_9(314) <= temp_mult_77(314);
partial_product_9(315) <= temp_mult_77(315);
partial_product_9(316) <= temp_mult_77(316);
partial_product_9(317) <= temp_mult_77(317);
partial_product_9(318) <= temp_mult_77(318);
partial_product_9(319) <= temp_mult_77(319);
partial_product_9(320) <= temp_mult_77(320);
partial_product_9(321) <= temp_mult_77(321);
partial_product_9(322) <= temp_mult_77(322);
partial_product_9(323) <= temp_mult_77(323);
partial_product_9(324) <= temp_mult_77(324);
partial_product_9(325) <= temp_mult_77(325);
partial_product_9(326) <= temp_mult_77(326);
partial_product_9(327) <= temp_mult_77(327);
partial_product_9(328) <= temp_mult_77(328);
partial_product_9(329) <= temp_mult_77(329);
partial_product_9(330) <= temp_mult_77(330);
partial_product_9(331) <= temp_mult_77(331);
partial_product_9(332) <= temp_mult_77(332);
partial_product_9(333) <= temp_mult_77(333);
partial_product_9(334) <= temp_mult_77(334);
partial_product_9(335) <= temp_mult_77(335);
partial_product_9(336) <= temp_mult_77(336);
partial_product_9(337) <= temp_mult_77(337);
partial_product_9(338) <= temp_mult_77(338);
partial_product_9(339) <= temp_mult_77(339);
partial_product_9(340) <= temp_mult_77(340);
partial_product_9(341) <= temp_mult_77(341);
partial_product_9(342) <= '0';
partial_product_9(343) <= '0';
partial_product_9(344) <= '0';
partial_product_9(345) <= '0';
partial_product_9(346) <= '0';
partial_product_9(347) <= '0';
partial_product_9(348) <= temp_mult_141(348);
partial_product_9(349) <= temp_mult_141(349);
partial_product_9(350) <= temp_mult_141(350);
partial_product_9(351) <= temp_mult_141(351);
partial_product_9(352) <= temp_mult_141(352);
partial_product_9(353) <= temp_mult_141(353);
partial_product_9(354) <= temp_mult_141(354);
partial_product_9(355) <= temp_mult_141(355);
partial_product_9(356) <= temp_mult_141(356);
partial_product_9(357) <= temp_mult_141(357);
partial_product_9(358) <= temp_mult_141(358);
partial_product_9(359) <= temp_mult_141(359);
partial_product_9(360) <= temp_mult_141(360);
partial_product_9(361) <= temp_mult_141(361);
partial_product_9(362) <= temp_mult_141(362);
partial_product_9(363) <= temp_mult_141(363);
partial_product_9(364) <= temp_mult_141(364);
partial_product_9(365) <= temp_mult_141(365);
partial_product_9(366) <= temp_mult_141(366);
partial_product_9(367) <= temp_mult_141(367);
partial_product_9(368) <= temp_mult_141(368);
partial_product_9(369) <= temp_mult_141(369);
partial_product_9(370) <= temp_mult_141(370);
partial_product_9(371) <= temp_mult_141(371);
partial_product_9(372) <= temp_mult_141(372);
partial_product_9(373) <= temp_mult_141(373);
partial_product_9(374) <= temp_mult_141(374);
partial_product_9(375) <= temp_mult_141(375);
partial_product_9(376) <= temp_mult_141(376);
partial_product_9(377) <= temp_mult_141(377);
partial_product_9(378) <= temp_mult_141(378);
partial_product_9(379) <= temp_mult_141(379);
partial_product_9(380) <= temp_mult_141(380);
partial_product_9(381) <= temp_mult_141(381);
partial_product_9(382) <= temp_mult_141(382);
partial_product_9(383) <= temp_mult_141(383);
partial_product_9(384) <= temp_mult_141(384);
partial_product_9(385) <= temp_mult_141(385);
partial_product_9(386) <= temp_mult_141(386);
partial_product_9(387) <= temp_mult_141(387);
partial_product_9(388) <= temp_mult_141(388);
partial_product_9(389) <= temp_mult_147(389);
partial_product_9(390) <= temp_mult_147(390);
partial_product_9(391) <= temp_mult_147(391);
partial_product_9(392) <= temp_mult_147(392);
partial_product_9(393) <= temp_mult_147(393);
partial_product_9(394) <= temp_mult_147(394);
partial_product_9(395) <= temp_mult_147(395);
partial_product_9(396) <= temp_mult_147(396);
partial_product_9(397) <= temp_mult_147(397);
partial_product_9(398) <= temp_mult_147(398);
partial_product_9(399) <= temp_mult_147(399);
partial_product_9(400) <= temp_mult_147(400);
partial_product_9(401) <= temp_mult_147(401);
partial_product_9(402) <= temp_mult_147(402);
partial_product_9(403) <= temp_mult_147(403);
partial_product_9(404) <= temp_mult_147(404);
partial_product_9(405) <= temp_mult_147(405);
partial_product_9(406) <= temp_mult_147(406);
partial_product_9(407) <= temp_mult_147(407);
partial_product_9(408) <= temp_mult_147(408);
partial_product_9(409) <= temp_mult_147(409);
partial_product_9(410) <= temp_mult_147(410);
partial_product_9(411) <= temp_mult_147(411);
partial_product_9(412) <= temp_mult_147(412);
partial_product_9(413) <= temp_mult_147(413);
partial_product_9(414) <= temp_mult_147(414);
partial_product_9(415) <= temp_mult_147(415);
partial_product_9(416) <= temp_mult_147(416);
partial_product_9(417) <= temp_mult_147(417);
partial_product_9(418) <= temp_mult_147(418);
partial_product_9(419) <= temp_mult_147(419);
partial_product_9(420) <= temp_mult_147(420);
partial_product_9(421) <= temp_mult_147(421);
partial_product_9(422) <= temp_mult_147(422);
partial_product_9(423) <= temp_mult_147(423);
partial_product_9(424) <= temp_mult_147(424);
partial_product_9(425) <= temp_mult_147(425);
partial_product_9(426) <= temp_mult_147(426);
partial_product_9(427) <= temp_mult_147(427);
partial_product_9(428) <= temp_mult_147(428);
partial_product_9(429) <= temp_mult_147(429);
partial_product_9(430) <= '0';
partial_product_9(431) <= '0';
partial_product_9(432) <= '0';
partial_product_9(433) <= '0';
partial_product_9(434) <= '0';
partial_product_9(435) <= '0';
partial_product_9(436) <= '0';
partial_product_9(437) <= '0';
partial_product_9(438) <= '0';
partial_product_9(439) <= '0';
partial_product_9(440) <= '0';
partial_product_9(441) <= '0';
partial_product_9(442) <= '0';
partial_product_9(443) <= '0';
partial_product_9(444) <= '0';
partial_product_9(445) <= '0';
partial_product_9(446) <= '0';
partial_product_9(447) <= '0';
partial_product_9(448) <= '0';
partial_product_9(449) <= '0';
partial_product_9(450) <= '0';
partial_product_9(451) <= '0';
partial_product_9(452) <= '0';
partial_product_9(453) <= '0';
partial_product_9(454) <= '0';
partial_product_9(455) <= '0';
partial_product_9(456) <= '0';
partial_product_9(457) <= '0';
partial_product_9(458) <= '0';
partial_product_9(459) <= '0';
partial_product_9(460) <= '0';
partial_product_9(461) <= '0';
partial_product_9(462) <= '0';
partial_product_9(463) <= '0';
partial_product_9(464) <= '0';
partial_product_9(465) <= '0';
partial_product_9(466) <= '0';
partial_product_9(467) <= '0';
partial_product_9(468) <= '0';
partial_product_9(469) <= '0';
partial_product_9(470) <= '0';
partial_product_9(471) <= '0';
partial_product_9(472) <= '0';
partial_product_9(473) <= '0';
partial_product_9(474) <= '0';
partial_product_9(475) <= '0';
partial_product_9(476) <= '0';
partial_product_9(477) <= '0';
partial_product_9(478) <= '0';
partial_product_9(479) <= '0';
partial_product_9(480) <= '0';
partial_product_9(481) <= '0';
partial_product_9(482) <= '0';
partial_product_9(483) <= '0';
partial_product_9(484) <= '0';
partial_product_9(485) <= '0';
partial_product_9(486) <= '0';
partial_product_9(487) <= '0';
partial_product_9(488) <= '0';
partial_product_9(489) <= '0';
partial_product_9(490) <= '0';
partial_product_9(491) <= '0';
partial_product_9(492) <= '0';
partial_product_9(493) <= '0';
partial_product_9(494) <= '0';
partial_product_9(495) <= '0';
partial_product_9(496) <= '0';
partial_product_9(497) <= '0';
partial_product_9(498) <= '0';
partial_product_9(499) <= '0';
partial_product_9(500) <= '0';
partial_product_9(501) <= '0';
partial_product_9(502) <= '0';
partial_product_9(503) <= '0';
partial_product_9(504) <= '0';
partial_product_9(505) <= '0';
partial_product_9(506) <= '0';
partial_product_9(507) <= '0';
partial_product_9(508) <= '0';
partial_product_9(509) <= '0';
partial_product_9(510) <= '0';
partial_product_9(511) <= '0';
partial_product_9(512) <= '0';
partial_product_10(0) <= '0';
partial_product_10(1) <= '0';
partial_product_10(2) <= '0';
partial_product_10(3) <= '0';
partial_product_10(4) <= '0';
partial_product_10(5) <= '0';
partial_product_10(6) <= '0';
partial_product_10(7) <= '0';
partial_product_10(8) <= '0';
partial_product_10(9) <= '0';
partial_product_10(10) <= '0';
partial_product_10(11) <= '0';
partial_product_10(12) <= '0';
partial_product_10(13) <= '0';
partial_product_10(14) <= '0';
partial_product_10(15) <= '0';
partial_product_10(16) <= '0';
partial_product_10(17) <= '0';
partial_product_10(18) <= '0';
partial_product_10(19) <= '0';
partial_product_10(20) <= '0';
partial_product_10(21) <= '0';
partial_product_10(22) <= '0';
partial_product_10(23) <= '0';
partial_product_10(24) <= '0';
partial_product_10(25) <= '0';
partial_product_10(26) <= '0';
partial_product_10(27) <= '0';
partial_product_10(28) <= '0';
partial_product_10(29) <= '0';
partial_product_10(30) <= '0';
partial_product_10(31) <= '0';
partial_product_10(32) <= '0';
partial_product_10(33) <= '0';
partial_product_10(34) <= '0';
partial_product_10(35) <= '0';
partial_product_10(36) <= '0';
partial_product_10(37) <= '0';
partial_product_10(38) <= '0';
partial_product_10(39) <= '0';
partial_product_10(40) <= '0';
partial_product_10(41) <= '0';
partial_product_10(42) <= '0';
partial_product_10(43) <= '0';
partial_product_10(44) <= '0';
partial_product_10(45) <= '0';
partial_product_10(46) <= '0';
partial_product_10(47) <= '0';
partial_product_10(48) <= '0';
partial_product_10(49) <= '0';
partial_product_10(50) <= '0';
partial_product_10(51) <= '0';
partial_product_10(52) <= '0';
partial_product_10(53) <= '0';
partial_product_10(54) <= '0';
partial_product_10(55) <= '0';
partial_product_10(56) <= '0';
partial_product_10(57) <= '0';
partial_product_10(58) <= '0';
partial_product_10(59) <= '0';
partial_product_10(60) <= '0';
partial_product_10(61) <= '0';
partial_product_10(62) <= '0';
partial_product_10(63) <= '0';
partial_product_10(64) <= '0';
partial_product_10(65) <= '0';
partial_product_10(66) <= '0';
partial_product_10(67) <= '0';
partial_product_10(68) <= '0';
partial_product_10(69) <= '0';
partial_product_10(70) <= '0';
partial_product_10(71) <= '0';
partial_product_10(72) <= '0';
partial_product_10(73) <= '0';
partial_product_10(74) <= '0';
partial_product_10(75) <= '0';
partial_product_10(76) <= '0';
partial_product_10(77) <= '0';
partial_product_10(78) <= '0';
partial_product_10(79) <= '0';
partial_product_10(80) <= '0';
partial_product_10(81) <= '0';
partial_product_10(82) <= '0';
partial_product_10(83) <= '0';
partial_product_10(84) <= '0';
partial_product_10(85) <= '0';
partial_product_10(86) <= '0';
partial_product_10(87) <= '0';
partial_product_10(88) <= '0';
partial_product_10(89) <= '0';
partial_product_10(90) <= '0';
partial_product_10(91) <= '0';
partial_product_10(92) <= '0';
partial_product_10(93) <= '0';
partial_product_10(94) <= '0';
partial_product_10(95) <= '0';
partial_product_10(96) <= '0';
partial_product_10(97) <= '0';
partial_product_10(98) <= '0';
partial_product_10(99) <= '0';
partial_product_10(100) <= '0';
partial_product_10(101) <= '0';
partial_product_10(102) <= temp_mult_30(102);
partial_product_10(103) <= temp_mult_30(103);
partial_product_10(104) <= temp_mult_30(104);
partial_product_10(105) <= temp_mult_30(105);
partial_product_10(106) <= temp_mult_30(106);
partial_product_10(107) <= temp_mult_30(107);
partial_product_10(108) <= temp_mult_30(108);
partial_product_10(109) <= temp_mult_30(109);
partial_product_10(110) <= temp_mult_30(110);
partial_product_10(111) <= temp_mult_30(111);
partial_product_10(112) <= temp_mult_30(112);
partial_product_10(113) <= temp_mult_30(113);
partial_product_10(114) <= temp_mult_30(114);
partial_product_10(115) <= temp_mult_30(115);
partial_product_10(116) <= temp_mult_30(116);
partial_product_10(117) <= temp_mult_30(117);
partial_product_10(118) <= temp_mult_30(118);
partial_product_10(119) <= temp_mult_30(119);
partial_product_10(120) <= temp_mult_30(120);
partial_product_10(121) <= temp_mult_30(121);
partial_product_10(122) <= temp_mult_30(122);
partial_product_10(123) <= temp_mult_30(123);
partial_product_10(124) <= temp_mult_30(124);
partial_product_10(125) <= temp_mult_30(125);
partial_product_10(126) <= temp_mult_30(126);
partial_product_10(127) <= temp_mult_30(127);
partial_product_10(128) <= temp_mult_30(128);
partial_product_10(129) <= temp_mult_30(129);
partial_product_10(130) <= temp_mult_30(130);
partial_product_10(131) <= temp_mult_30(131);
partial_product_10(132) <= temp_mult_30(132);
partial_product_10(133) <= temp_mult_30(133);
partial_product_10(134) <= temp_mult_30(134);
partial_product_10(135) <= temp_mult_30(135);
partial_product_10(136) <= temp_mult_30(136);
partial_product_10(137) <= temp_mult_30(137);
partial_product_10(138) <= temp_mult_30(138);
partial_product_10(139) <= temp_mult_30(139);
partial_product_10(140) <= temp_mult_30(140);
partial_product_10(141) <= temp_mult_30(141);
partial_product_10(142) <= temp_mult_30(142);
partial_product_10(143) <= temp_mult_36(143);
partial_product_10(144) <= temp_mult_36(144);
partial_product_10(145) <= temp_mult_36(145);
partial_product_10(146) <= temp_mult_36(146);
partial_product_10(147) <= temp_mult_36(147);
partial_product_10(148) <= temp_mult_36(148);
partial_product_10(149) <= temp_mult_36(149);
partial_product_10(150) <= temp_mult_36(150);
partial_product_10(151) <= temp_mult_36(151);
partial_product_10(152) <= temp_mult_36(152);
partial_product_10(153) <= temp_mult_36(153);
partial_product_10(154) <= temp_mult_36(154);
partial_product_10(155) <= temp_mult_36(155);
partial_product_10(156) <= temp_mult_36(156);
partial_product_10(157) <= temp_mult_36(157);
partial_product_10(158) <= temp_mult_36(158);
partial_product_10(159) <= temp_mult_36(159);
partial_product_10(160) <= temp_mult_36(160);
partial_product_10(161) <= temp_mult_36(161);
partial_product_10(162) <= temp_mult_36(162);
partial_product_10(163) <= temp_mult_36(163);
partial_product_10(164) <= temp_mult_36(164);
partial_product_10(165) <= temp_mult_36(165);
partial_product_10(166) <= temp_mult_36(166);
partial_product_10(167) <= temp_mult_36(167);
partial_product_10(168) <= temp_mult_36(168);
partial_product_10(169) <= temp_mult_36(169);
partial_product_10(170) <= temp_mult_36(170);
partial_product_10(171) <= temp_mult_36(171);
partial_product_10(172) <= temp_mult_36(172);
partial_product_10(173) <= temp_mult_36(173);
partial_product_10(174) <= temp_mult_36(174);
partial_product_10(175) <= temp_mult_36(175);
partial_product_10(176) <= temp_mult_36(176);
partial_product_10(177) <= temp_mult_36(177);
partial_product_10(178) <= temp_mult_36(178);
partial_product_10(179) <= temp_mult_36(179);
partial_product_10(180) <= temp_mult_36(180);
partial_product_10(181) <= temp_mult_36(181);
partial_product_10(182) <= temp_mult_36(182);
partial_product_10(183) <= temp_mult_36(183);
partial_product_10(184) <= temp_mult_96(184);
partial_product_10(185) <= temp_mult_96(185);
partial_product_10(186) <= temp_mult_96(186);
partial_product_10(187) <= temp_mult_96(187);
partial_product_10(188) <= temp_mult_96(188);
partial_product_10(189) <= temp_mult_96(189);
partial_product_10(190) <= temp_mult_96(190);
partial_product_10(191) <= temp_mult_96(191);
partial_product_10(192) <= temp_mult_96(192);
partial_product_10(193) <= temp_mult_96(193);
partial_product_10(194) <= temp_mult_96(194);
partial_product_10(195) <= temp_mult_96(195);
partial_product_10(196) <= temp_mult_96(196);
partial_product_10(197) <= temp_mult_96(197);
partial_product_10(198) <= temp_mult_96(198);
partial_product_10(199) <= temp_mult_96(199);
partial_product_10(200) <= temp_mult_96(200);
partial_product_10(201) <= temp_mult_96(201);
partial_product_10(202) <= temp_mult_96(202);
partial_product_10(203) <= temp_mult_96(203);
partial_product_10(204) <= temp_mult_96(204);
partial_product_10(205) <= temp_mult_96(205);
partial_product_10(206) <= temp_mult_96(206);
partial_product_10(207) <= temp_mult_96(207);
partial_product_10(208) <= temp_mult_96(208);
partial_product_10(209) <= temp_mult_96(209);
partial_product_10(210) <= temp_mult_96(210);
partial_product_10(211) <= temp_mult_96(211);
partial_product_10(212) <= temp_mult_96(212);
partial_product_10(213) <= temp_mult_96(213);
partial_product_10(214) <= temp_mult_96(214);
partial_product_10(215) <= temp_mult_96(215);
partial_product_10(216) <= temp_mult_96(216);
partial_product_10(217) <= temp_mult_96(217);
partial_product_10(218) <= temp_mult_96(218);
partial_product_10(219) <= temp_mult_96(219);
partial_product_10(220) <= temp_mult_96(220);
partial_product_10(221) <= temp_mult_96(221);
partial_product_10(222) <= temp_mult_96(222);
partial_product_10(223) <= temp_mult_96(223);
partial_product_10(224) <= temp_mult_96(224);
partial_product_10(225) <= temp_mult_105(225);
partial_product_10(226) <= temp_mult_105(226);
partial_product_10(227) <= temp_mult_105(227);
partial_product_10(228) <= temp_mult_105(228);
partial_product_10(229) <= temp_mult_105(229);
partial_product_10(230) <= temp_mult_105(230);
partial_product_10(231) <= temp_mult_105(231);
partial_product_10(232) <= temp_mult_105(232);
partial_product_10(233) <= temp_mult_105(233);
partial_product_10(234) <= temp_mult_105(234);
partial_product_10(235) <= temp_mult_105(235);
partial_product_10(236) <= temp_mult_105(236);
partial_product_10(237) <= temp_mult_105(237);
partial_product_10(238) <= temp_mult_105(238);
partial_product_10(239) <= temp_mult_105(239);
partial_product_10(240) <= temp_mult_105(240);
partial_product_10(241) <= temp_mult_105(241);
partial_product_10(242) <= temp_mult_105(242);
partial_product_10(243) <= temp_mult_105(243);
partial_product_10(244) <= temp_mult_105(244);
partial_product_10(245) <= temp_mult_105(245);
partial_product_10(246) <= temp_mult_105(246);
partial_product_10(247) <= temp_mult_105(247);
partial_product_10(248) <= temp_mult_105(248);
partial_product_10(249) <= temp_mult_105(249);
partial_product_10(250) <= temp_mult_105(250);
partial_product_10(251) <= temp_mult_105(251);
partial_product_10(252) <= temp_mult_105(252);
partial_product_10(253) <= temp_mult_105(253);
partial_product_10(254) <= temp_mult_105(254);
partial_product_10(255) <= temp_mult_105(255);
partial_product_10(256) <= temp_mult_105(256);
partial_product_10(257) <= temp_mult_105(257);
partial_product_10(258) <= temp_mult_105(258);
partial_product_10(259) <= temp_mult_105(259);
partial_product_10(260) <= temp_mult_105(260);
partial_product_10(261) <= temp_mult_105(261);
partial_product_10(262) <= temp_mult_105(262);
partial_product_10(263) <= temp_mult_105(263);
partial_product_10(264) <= temp_mult_105(264);
partial_product_10(265) <= temp_mult_105(265);
partial_product_10(266) <= temp_mult_114(266);
partial_product_10(267) <= temp_mult_114(267);
partial_product_10(268) <= temp_mult_114(268);
partial_product_10(269) <= temp_mult_114(269);
partial_product_10(270) <= temp_mult_114(270);
partial_product_10(271) <= temp_mult_114(271);
partial_product_10(272) <= temp_mult_114(272);
partial_product_10(273) <= temp_mult_114(273);
partial_product_10(274) <= temp_mult_114(274);
partial_product_10(275) <= temp_mult_114(275);
partial_product_10(276) <= temp_mult_114(276);
partial_product_10(277) <= temp_mult_114(277);
partial_product_10(278) <= temp_mult_114(278);
partial_product_10(279) <= temp_mult_114(279);
partial_product_10(280) <= temp_mult_114(280);
partial_product_10(281) <= temp_mult_114(281);
partial_product_10(282) <= temp_mult_114(282);
partial_product_10(283) <= temp_mult_114(283);
partial_product_10(284) <= temp_mult_114(284);
partial_product_10(285) <= temp_mult_114(285);
partial_product_10(286) <= temp_mult_114(286);
partial_product_10(287) <= temp_mult_114(287);
partial_product_10(288) <= temp_mult_114(288);
partial_product_10(289) <= temp_mult_114(289);
partial_product_10(290) <= temp_mult_114(290);
partial_product_10(291) <= temp_mult_114(291);
partial_product_10(292) <= temp_mult_114(292);
partial_product_10(293) <= temp_mult_114(293);
partial_product_10(294) <= temp_mult_114(294);
partial_product_10(295) <= temp_mult_114(295);
partial_product_10(296) <= temp_mult_114(296);
partial_product_10(297) <= temp_mult_114(297);
partial_product_10(298) <= temp_mult_114(298);
partial_product_10(299) <= temp_mult_114(299);
partial_product_10(300) <= temp_mult_114(300);
partial_product_10(301) <= temp_mult_114(301);
partial_product_10(302) <= temp_mult_114(302);
partial_product_10(303) <= temp_mult_114(303);
partial_product_10(304) <= temp_mult_114(304);
partial_product_10(305) <= temp_mult_114(305);
partial_product_10(306) <= temp_mult_114(306);
partial_product_10(307) <= temp_mult_135(307);
partial_product_10(308) <= temp_mult_135(308);
partial_product_10(309) <= temp_mult_135(309);
partial_product_10(310) <= temp_mult_135(310);
partial_product_10(311) <= temp_mult_135(311);
partial_product_10(312) <= temp_mult_135(312);
partial_product_10(313) <= temp_mult_135(313);
partial_product_10(314) <= temp_mult_135(314);
partial_product_10(315) <= temp_mult_135(315);
partial_product_10(316) <= temp_mult_135(316);
partial_product_10(317) <= temp_mult_135(317);
partial_product_10(318) <= temp_mult_135(318);
partial_product_10(319) <= temp_mult_135(319);
partial_product_10(320) <= temp_mult_135(320);
partial_product_10(321) <= temp_mult_135(321);
partial_product_10(322) <= temp_mult_135(322);
partial_product_10(323) <= temp_mult_135(323);
partial_product_10(324) <= temp_mult_135(324);
partial_product_10(325) <= temp_mult_135(325);
partial_product_10(326) <= temp_mult_135(326);
partial_product_10(327) <= temp_mult_135(327);
partial_product_10(328) <= temp_mult_135(328);
partial_product_10(329) <= temp_mult_135(329);
partial_product_10(330) <= temp_mult_135(330);
partial_product_10(331) <= temp_mult_135(331);
partial_product_10(332) <= temp_mult_135(332);
partial_product_10(333) <= temp_mult_135(333);
partial_product_10(334) <= temp_mult_135(334);
partial_product_10(335) <= temp_mult_135(335);
partial_product_10(336) <= temp_mult_135(336);
partial_product_10(337) <= temp_mult_135(337);
partial_product_10(338) <= temp_mult_135(338);
partial_product_10(339) <= temp_mult_135(339);
partial_product_10(340) <= temp_mult_135(340);
partial_product_10(341) <= temp_mult_135(341);
partial_product_10(342) <= temp_mult_135(342);
partial_product_10(343) <= temp_mult_135(343);
partial_product_10(344) <= temp_mult_135(344);
partial_product_10(345) <= temp_mult_135(345);
partial_product_10(346) <= temp_mult_135(346);
partial_product_10(347) <= temp_mult_135(347);
partial_product_10(348) <= '0';
partial_product_10(349) <= '0';
partial_product_10(350) <= '0';
partial_product_10(351) <= temp_mult_119(351);
partial_product_10(352) <= temp_mult_119(352);
partial_product_10(353) <= temp_mult_119(353);
partial_product_10(354) <= temp_mult_119(354);
partial_product_10(355) <= temp_mult_119(355);
partial_product_10(356) <= temp_mult_119(356);
partial_product_10(357) <= temp_mult_119(357);
partial_product_10(358) <= temp_mult_119(358);
partial_product_10(359) <= temp_mult_119(359);
partial_product_10(360) <= temp_mult_119(360);
partial_product_10(361) <= temp_mult_119(361);
partial_product_10(362) <= temp_mult_119(362);
partial_product_10(363) <= temp_mult_119(363);
partial_product_10(364) <= temp_mult_119(364);
partial_product_10(365) <= temp_mult_119(365);
partial_product_10(366) <= temp_mult_119(366);
partial_product_10(367) <= temp_mult_119(367);
partial_product_10(368) <= temp_mult_119(368);
partial_product_10(369) <= temp_mult_119(369);
partial_product_10(370) <= temp_mult_119(370);
partial_product_10(371) <= temp_mult_119(371);
partial_product_10(372) <= temp_mult_119(372);
partial_product_10(373) <= temp_mult_119(373);
partial_product_10(374) <= temp_mult_119(374);
partial_product_10(375) <= temp_mult_119(375);
partial_product_10(376) <= temp_mult_119(376);
partial_product_10(377) <= temp_mult_119(377);
partial_product_10(378) <= temp_mult_119(378);
partial_product_10(379) <= temp_mult_119(379);
partial_product_10(380) <= temp_mult_119(380);
partial_product_10(381) <= temp_mult_119(381);
partial_product_10(382) <= temp_mult_119(382);
partial_product_10(383) <= temp_mult_119(383);
partial_product_10(384) <= temp_mult_119(384);
partial_product_10(385) <= temp_mult_119(385);
partial_product_10(386) <= temp_mult_119(386);
partial_product_10(387) <= temp_mult_119(387);
partial_product_10(388) <= temp_mult_119(388);
partial_product_10(389) <= temp_mult_119(389);
partial_product_10(390) <= temp_mult_119(390);
partial_product_10(391) <= temp_mult_119(391);
partial_product_10(392) <= '0';
partial_product_10(393) <= '0';
partial_product_10(394) <= '0';
partial_product_10(395) <= '0';
partial_product_10(396) <= '0';
partial_product_10(397) <= '0';
partial_product_10(398) <= '0';
partial_product_10(399) <= '0';
partial_product_10(400) <= '0';
partial_product_10(401) <= '0';
partial_product_10(402) <= '0';
partial_product_10(403) <= '0';
partial_product_10(404) <= '0';
partial_product_10(405) <= '0';
partial_product_10(406) <= '0';
partial_product_10(407) <= '0';
partial_product_10(408) <= '0';
partial_product_10(409) <= '0';
partial_product_10(410) <= '0';
partial_product_10(411) <= '0';
partial_product_10(412) <= '0';
partial_product_10(413) <= '0';
partial_product_10(414) <= '0';
partial_product_10(415) <= '0';
partial_product_10(416) <= '0';
partial_product_10(417) <= '0';
partial_product_10(418) <= '0';
partial_product_10(419) <= '0';
partial_product_10(420) <= '0';
partial_product_10(421) <= '0';
partial_product_10(422) <= '0';
partial_product_10(423) <= '0';
partial_product_10(424) <= '0';
partial_product_10(425) <= '0';
partial_product_10(426) <= '0';
partial_product_10(427) <= '0';
partial_product_10(428) <= '0';
partial_product_10(429) <= '0';
partial_product_10(430) <= '0';
partial_product_10(431) <= '0';
partial_product_10(432) <= '0';
partial_product_10(433) <= '0';
partial_product_10(434) <= '0';
partial_product_10(435) <= '0';
partial_product_10(436) <= '0';
partial_product_10(437) <= '0';
partial_product_10(438) <= '0';
partial_product_10(439) <= '0';
partial_product_10(440) <= '0';
partial_product_10(441) <= '0';
partial_product_10(442) <= '0';
partial_product_10(443) <= '0';
partial_product_10(444) <= '0';
partial_product_10(445) <= '0';
partial_product_10(446) <= '0';
partial_product_10(447) <= '0';
partial_product_10(448) <= '0';
partial_product_10(449) <= '0';
partial_product_10(450) <= '0';
partial_product_10(451) <= '0';
partial_product_10(452) <= '0';
partial_product_10(453) <= '0';
partial_product_10(454) <= '0';
partial_product_10(455) <= '0';
partial_product_10(456) <= '0';
partial_product_10(457) <= '0';
partial_product_10(458) <= '0';
partial_product_10(459) <= '0';
partial_product_10(460) <= '0';
partial_product_10(461) <= '0';
partial_product_10(462) <= '0';
partial_product_10(463) <= '0';
partial_product_10(464) <= '0';
partial_product_10(465) <= '0';
partial_product_10(466) <= '0';
partial_product_10(467) <= '0';
partial_product_10(468) <= '0';
partial_product_10(469) <= '0';
partial_product_10(470) <= '0';
partial_product_10(471) <= '0';
partial_product_10(472) <= '0';
partial_product_10(473) <= '0';
partial_product_10(474) <= '0';
partial_product_10(475) <= '0';
partial_product_10(476) <= '0';
partial_product_10(477) <= '0';
partial_product_10(478) <= '0';
partial_product_10(479) <= '0';
partial_product_10(480) <= '0';
partial_product_10(481) <= '0';
partial_product_10(482) <= '0';
partial_product_10(483) <= '0';
partial_product_10(484) <= '0';
partial_product_10(485) <= '0';
partial_product_10(486) <= '0';
partial_product_10(487) <= '0';
partial_product_10(488) <= '0';
partial_product_10(489) <= '0';
partial_product_10(490) <= '0';
partial_product_10(491) <= '0';
partial_product_10(492) <= '0';
partial_product_10(493) <= '0';
partial_product_10(494) <= '0';
partial_product_10(495) <= '0';
partial_product_10(496) <= '0';
partial_product_10(497) <= '0';
partial_product_10(498) <= '0';
partial_product_10(499) <= '0';
partial_product_10(500) <= '0';
partial_product_10(501) <= '0';
partial_product_10(502) <= '0';
partial_product_10(503) <= '0';
partial_product_10(504) <= '0';
partial_product_10(505) <= '0';
partial_product_10(506) <= '0';
partial_product_10(507) <= '0';
partial_product_10(508) <= '0';
partial_product_10(509) <= '0';
partial_product_10(510) <= '0';
partial_product_10(511) <= '0';
partial_product_10(512) <= '0';
partial_product_11(0) <= '0';
partial_product_11(1) <= '0';
partial_product_11(2) <= '0';
partial_product_11(3) <= '0';
partial_product_11(4) <= '0';
partial_product_11(5) <= '0';
partial_product_11(6) <= '0';
partial_product_11(7) <= '0';
partial_product_11(8) <= '0';
partial_product_11(9) <= '0';
partial_product_11(10) <= '0';
partial_product_11(11) <= '0';
partial_product_11(12) <= '0';
partial_product_11(13) <= '0';
partial_product_11(14) <= '0';
partial_product_11(15) <= '0';
partial_product_11(16) <= '0';
partial_product_11(17) <= '0';
partial_product_11(18) <= '0';
partial_product_11(19) <= '0';
partial_product_11(20) <= '0';
partial_product_11(21) <= '0';
partial_product_11(22) <= '0';
partial_product_11(23) <= '0';
partial_product_11(24) <= '0';
partial_product_11(25) <= '0';
partial_product_11(26) <= '0';
partial_product_11(27) <= '0';
partial_product_11(28) <= '0';
partial_product_11(29) <= '0';
partial_product_11(30) <= '0';
partial_product_11(31) <= '0';
partial_product_11(32) <= '0';
partial_product_11(33) <= '0';
partial_product_11(34) <= '0';
partial_product_11(35) <= '0';
partial_product_11(36) <= '0';
partial_product_11(37) <= '0';
partial_product_11(38) <= '0';
partial_product_11(39) <= '0';
partial_product_11(40) <= '0';
partial_product_11(41) <= '0';
partial_product_11(42) <= '0';
partial_product_11(43) <= '0';
partial_product_11(44) <= '0';
partial_product_11(45) <= '0';
partial_product_11(46) <= '0';
partial_product_11(47) <= '0';
partial_product_11(48) <= '0';
partial_product_11(49) <= '0';
partial_product_11(50) <= '0';
partial_product_11(51) <= '0';
partial_product_11(52) <= '0';
partial_product_11(53) <= '0';
partial_product_11(54) <= '0';
partial_product_11(55) <= '0';
partial_product_11(56) <= '0';
partial_product_11(57) <= '0';
partial_product_11(58) <= '0';
partial_product_11(59) <= '0';
partial_product_11(60) <= '0';
partial_product_11(61) <= '0';
partial_product_11(62) <= '0';
partial_product_11(63) <= '0';
partial_product_11(64) <= '0';
partial_product_11(65) <= '0';
partial_product_11(66) <= '0';
partial_product_11(67) <= '0';
partial_product_11(68) <= '0';
partial_product_11(69) <= '0';
partial_product_11(70) <= '0';
partial_product_11(71) <= '0';
partial_product_11(72) <= '0';
partial_product_11(73) <= '0';
partial_product_11(74) <= '0';
partial_product_11(75) <= '0';
partial_product_11(76) <= '0';
partial_product_11(77) <= '0';
partial_product_11(78) <= '0';
partial_product_11(79) <= '0';
partial_product_11(80) <= '0';
partial_product_11(81) <= '0';
partial_product_11(82) <= '0';
partial_product_11(83) <= '0';
partial_product_11(84) <= '0';
partial_product_11(85) <= '0';
partial_product_11(86) <= '0';
partial_product_11(87) <= '0';
partial_product_11(88) <= '0';
partial_product_11(89) <= '0';
partial_product_11(90) <= '0';
partial_product_11(91) <= '0';
partial_product_11(92) <= '0';
partial_product_11(93) <= '0';
partial_product_11(94) <= '0';
partial_product_11(95) <= '0';
partial_product_11(96) <= '0';
partial_product_11(97) <= '0';
partial_product_11(98) <= '0';
partial_product_11(99) <= '0';
partial_product_11(100) <= '0';
partial_product_11(101) <= '0';
partial_product_11(102) <= '0';
partial_product_11(103) <= '0';
partial_product_11(104) <= '0';
partial_product_11(105) <= '0';
partial_product_11(106) <= '0';
partial_product_11(107) <= '0';
partial_product_11(108) <= '0';
partial_product_11(109) <= '0';
partial_product_11(110) <= '0';
partial_product_11(111) <= '0';
partial_product_11(112) <= '0';
partial_product_11(113) <= '0';
partial_product_11(114) <= '0';
partial_product_11(115) <= '0';
partial_product_11(116) <= '0';
partial_product_11(117) <= '0';
partial_product_11(118) <= '0';
partial_product_11(119) <= temp_mult_35(119);
partial_product_11(120) <= temp_mult_35(120);
partial_product_11(121) <= temp_mult_35(121);
partial_product_11(122) <= temp_mult_35(122);
partial_product_11(123) <= temp_mult_35(123);
partial_product_11(124) <= temp_mult_35(124);
partial_product_11(125) <= temp_mult_35(125);
partial_product_11(126) <= temp_mult_35(126);
partial_product_11(127) <= temp_mult_35(127);
partial_product_11(128) <= temp_mult_35(128);
partial_product_11(129) <= temp_mult_35(129);
partial_product_11(130) <= temp_mult_35(130);
partial_product_11(131) <= temp_mult_35(131);
partial_product_11(132) <= temp_mult_35(132);
partial_product_11(133) <= temp_mult_35(133);
partial_product_11(134) <= temp_mult_35(134);
partial_product_11(135) <= temp_mult_35(135);
partial_product_11(136) <= temp_mult_35(136);
partial_product_11(137) <= temp_mult_35(137);
partial_product_11(138) <= temp_mult_35(138);
partial_product_11(139) <= temp_mult_35(139);
partial_product_11(140) <= temp_mult_35(140);
partial_product_11(141) <= temp_mult_35(141);
partial_product_11(142) <= temp_mult_35(142);
partial_product_11(143) <= temp_mult_35(143);
partial_product_11(144) <= temp_mult_35(144);
partial_product_11(145) <= temp_mult_35(145);
partial_product_11(146) <= temp_mult_35(146);
partial_product_11(147) <= temp_mult_35(147);
partial_product_11(148) <= temp_mult_35(148);
partial_product_11(149) <= temp_mult_35(149);
partial_product_11(150) <= temp_mult_35(150);
partial_product_11(151) <= temp_mult_35(151);
partial_product_11(152) <= temp_mult_35(152);
partial_product_11(153) <= temp_mult_35(153);
partial_product_11(154) <= temp_mult_35(154);
partial_product_11(155) <= temp_mult_35(155);
partial_product_11(156) <= temp_mult_35(156);
partial_product_11(157) <= temp_mult_35(157);
partial_product_11(158) <= temp_mult_35(158);
partial_product_11(159) <= temp_mult_35(159);
partial_product_11(160) <= temp_mult_88(160);
partial_product_11(161) <= temp_mult_88(161);
partial_product_11(162) <= temp_mult_88(162);
partial_product_11(163) <= temp_mult_88(163);
partial_product_11(164) <= temp_mult_88(164);
partial_product_11(165) <= temp_mult_88(165);
partial_product_11(166) <= temp_mult_88(166);
partial_product_11(167) <= temp_mult_88(167);
partial_product_11(168) <= temp_mult_88(168);
partial_product_11(169) <= temp_mult_88(169);
partial_product_11(170) <= temp_mult_88(170);
partial_product_11(171) <= temp_mult_88(171);
partial_product_11(172) <= temp_mult_88(172);
partial_product_11(173) <= temp_mult_88(173);
partial_product_11(174) <= temp_mult_88(174);
partial_product_11(175) <= temp_mult_88(175);
partial_product_11(176) <= temp_mult_88(176);
partial_product_11(177) <= temp_mult_88(177);
partial_product_11(178) <= temp_mult_88(178);
partial_product_11(179) <= temp_mult_88(179);
partial_product_11(180) <= temp_mult_88(180);
partial_product_11(181) <= temp_mult_88(181);
partial_product_11(182) <= temp_mult_88(182);
partial_product_11(183) <= temp_mult_88(183);
partial_product_11(184) <= temp_mult_88(184);
partial_product_11(185) <= temp_mult_88(185);
partial_product_11(186) <= temp_mult_88(186);
partial_product_11(187) <= temp_mult_88(187);
partial_product_11(188) <= temp_mult_88(188);
partial_product_11(189) <= temp_mult_88(189);
partial_product_11(190) <= temp_mult_88(190);
partial_product_11(191) <= temp_mult_88(191);
partial_product_11(192) <= temp_mult_88(192);
partial_product_11(193) <= temp_mult_88(193);
partial_product_11(194) <= temp_mult_88(194);
partial_product_11(195) <= temp_mult_88(195);
partial_product_11(196) <= temp_mult_88(196);
partial_product_11(197) <= temp_mult_88(197);
partial_product_11(198) <= temp_mult_88(198);
partial_product_11(199) <= temp_mult_88(199);
partial_product_11(200) <= temp_mult_88(200);
partial_product_11(201) <= temp_mult_97(201);
partial_product_11(202) <= temp_mult_97(202);
partial_product_11(203) <= temp_mult_97(203);
partial_product_11(204) <= temp_mult_97(204);
partial_product_11(205) <= temp_mult_97(205);
partial_product_11(206) <= temp_mult_97(206);
partial_product_11(207) <= temp_mult_97(207);
partial_product_11(208) <= temp_mult_97(208);
partial_product_11(209) <= temp_mult_97(209);
partial_product_11(210) <= temp_mult_97(210);
partial_product_11(211) <= temp_mult_97(211);
partial_product_11(212) <= temp_mult_97(212);
partial_product_11(213) <= temp_mult_97(213);
partial_product_11(214) <= temp_mult_97(214);
partial_product_11(215) <= temp_mult_97(215);
partial_product_11(216) <= temp_mult_97(216);
partial_product_11(217) <= temp_mult_97(217);
partial_product_11(218) <= temp_mult_97(218);
partial_product_11(219) <= temp_mult_97(219);
partial_product_11(220) <= temp_mult_97(220);
partial_product_11(221) <= temp_mult_97(221);
partial_product_11(222) <= temp_mult_97(222);
partial_product_11(223) <= temp_mult_97(223);
partial_product_11(224) <= temp_mult_97(224);
partial_product_11(225) <= temp_mult_97(225);
partial_product_11(226) <= temp_mult_97(226);
partial_product_11(227) <= temp_mult_97(227);
partial_product_11(228) <= temp_mult_97(228);
partial_product_11(229) <= temp_mult_97(229);
partial_product_11(230) <= temp_mult_97(230);
partial_product_11(231) <= temp_mult_97(231);
partial_product_11(232) <= temp_mult_97(232);
partial_product_11(233) <= temp_mult_97(233);
partial_product_11(234) <= temp_mult_97(234);
partial_product_11(235) <= temp_mult_97(235);
partial_product_11(236) <= temp_mult_97(236);
partial_product_11(237) <= temp_mult_97(237);
partial_product_11(238) <= temp_mult_97(238);
partial_product_11(239) <= temp_mult_97(239);
partial_product_11(240) <= temp_mult_97(240);
partial_product_11(241) <= temp_mult_97(241);
partial_product_11(242) <= temp_mult_106(242);
partial_product_11(243) <= temp_mult_106(243);
partial_product_11(244) <= temp_mult_106(244);
partial_product_11(245) <= temp_mult_106(245);
partial_product_11(246) <= temp_mult_106(246);
partial_product_11(247) <= temp_mult_106(247);
partial_product_11(248) <= temp_mult_106(248);
partial_product_11(249) <= temp_mult_106(249);
partial_product_11(250) <= temp_mult_106(250);
partial_product_11(251) <= temp_mult_106(251);
partial_product_11(252) <= temp_mult_106(252);
partial_product_11(253) <= temp_mult_106(253);
partial_product_11(254) <= temp_mult_106(254);
partial_product_11(255) <= temp_mult_106(255);
partial_product_11(256) <= temp_mult_106(256);
partial_product_11(257) <= temp_mult_106(257);
partial_product_11(258) <= temp_mult_106(258);
partial_product_11(259) <= temp_mult_106(259);
partial_product_11(260) <= temp_mult_106(260);
partial_product_11(261) <= temp_mult_106(261);
partial_product_11(262) <= temp_mult_106(262);
partial_product_11(263) <= temp_mult_106(263);
partial_product_11(264) <= temp_mult_106(264);
partial_product_11(265) <= temp_mult_106(265);
partial_product_11(266) <= temp_mult_106(266);
partial_product_11(267) <= temp_mult_106(267);
partial_product_11(268) <= temp_mult_106(268);
partial_product_11(269) <= temp_mult_106(269);
partial_product_11(270) <= temp_mult_106(270);
partial_product_11(271) <= temp_mult_106(271);
partial_product_11(272) <= temp_mult_106(272);
partial_product_11(273) <= temp_mult_106(273);
partial_product_11(274) <= temp_mult_106(274);
partial_product_11(275) <= temp_mult_106(275);
partial_product_11(276) <= temp_mult_106(276);
partial_product_11(277) <= temp_mult_106(277);
partial_product_11(278) <= temp_mult_106(278);
partial_product_11(279) <= temp_mult_106(279);
partial_product_11(280) <= temp_mult_106(280);
partial_product_11(281) <= temp_mult_106(281);
partial_product_11(282) <= temp_mult_106(282);
partial_product_11(283) <= temp_mult_115(283);
partial_product_11(284) <= temp_mult_115(284);
partial_product_11(285) <= temp_mult_115(285);
partial_product_11(286) <= temp_mult_115(286);
partial_product_11(287) <= temp_mult_115(287);
partial_product_11(288) <= temp_mult_115(288);
partial_product_11(289) <= temp_mult_115(289);
partial_product_11(290) <= temp_mult_115(290);
partial_product_11(291) <= temp_mult_115(291);
partial_product_11(292) <= temp_mult_115(292);
partial_product_11(293) <= temp_mult_115(293);
partial_product_11(294) <= temp_mult_115(294);
partial_product_11(295) <= temp_mult_115(295);
partial_product_11(296) <= temp_mult_115(296);
partial_product_11(297) <= temp_mult_115(297);
partial_product_11(298) <= temp_mult_115(298);
partial_product_11(299) <= temp_mult_115(299);
partial_product_11(300) <= temp_mult_115(300);
partial_product_11(301) <= temp_mult_115(301);
partial_product_11(302) <= temp_mult_115(302);
partial_product_11(303) <= temp_mult_115(303);
partial_product_11(304) <= temp_mult_115(304);
partial_product_11(305) <= temp_mult_115(305);
partial_product_11(306) <= temp_mult_115(306);
partial_product_11(307) <= temp_mult_115(307);
partial_product_11(308) <= temp_mult_115(308);
partial_product_11(309) <= temp_mult_115(309);
partial_product_11(310) <= temp_mult_115(310);
partial_product_11(311) <= temp_mult_115(311);
partial_product_11(312) <= temp_mult_115(312);
partial_product_11(313) <= temp_mult_115(313);
partial_product_11(314) <= temp_mult_115(314);
partial_product_11(315) <= temp_mult_115(315);
partial_product_11(316) <= temp_mult_115(316);
partial_product_11(317) <= temp_mult_115(317);
partial_product_11(318) <= temp_mult_115(318);
partial_product_11(319) <= temp_mult_115(319);
partial_product_11(320) <= temp_mult_115(320);
partial_product_11(321) <= temp_mult_115(321);
partial_product_11(322) <= temp_mult_115(322);
partial_product_11(323) <= temp_mult_115(323);
partial_product_11(324) <= temp_mult_140(324);
partial_product_11(325) <= temp_mult_140(325);
partial_product_11(326) <= temp_mult_140(326);
partial_product_11(327) <= temp_mult_140(327);
partial_product_11(328) <= temp_mult_140(328);
partial_product_11(329) <= temp_mult_140(329);
partial_product_11(330) <= temp_mult_140(330);
partial_product_11(331) <= temp_mult_140(331);
partial_product_11(332) <= temp_mult_140(332);
partial_product_11(333) <= temp_mult_140(333);
partial_product_11(334) <= temp_mult_140(334);
partial_product_11(335) <= temp_mult_140(335);
partial_product_11(336) <= temp_mult_140(336);
partial_product_11(337) <= temp_mult_140(337);
partial_product_11(338) <= temp_mult_140(338);
partial_product_11(339) <= temp_mult_140(339);
partial_product_11(340) <= temp_mult_140(340);
partial_product_11(341) <= temp_mult_140(341);
partial_product_11(342) <= temp_mult_140(342);
partial_product_11(343) <= temp_mult_140(343);
partial_product_11(344) <= temp_mult_140(344);
partial_product_11(345) <= temp_mult_140(345);
partial_product_11(346) <= temp_mult_140(346);
partial_product_11(347) <= temp_mult_140(347);
partial_product_11(348) <= temp_mult_140(348);
partial_product_11(349) <= temp_mult_140(349);
partial_product_11(350) <= temp_mult_140(350);
partial_product_11(351) <= temp_mult_140(351);
partial_product_11(352) <= temp_mult_140(352);
partial_product_11(353) <= temp_mult_140(353);
partial_product_11(354) <= temp_mult_140(354);
partial_product_11(355) <= temp_mult_140(355);
partial_product_11(356) <= temp_mult_140(356);
partial_product_11(357) <= temp_mult_140(357);
partial_product_11(358) <= temp_mult_140(358);
partial_product_11(359) <= temp_mult_140(359);
partial_product_11(360) <= temp_mult_140(360);
partial_product_11(361) <= temp_mult_140(361);
partial_product_11(362) <= temp_mult_140(362);
partial_product_11(363) <= temp_mult_140(363);
partial_product_11(364) <= temp_mult_140(364);
partial_product_11(365) <= '0';
partial_product_11(366) <= '0';
partial_product_11(367) <= '0';
partial_product_11(368) <= '0';
partial_product_11(369) <= '0';
partial_product_11(370) <= '0';
partial_product_11(371) <= '0';
partial_product_11(372) <= '0';
partial_product_11(373) <= '0';
partial_product_11(374) <= '0';
partial_product_11(375) <= temp_mult_155(375);
partial_product_11(376) <= temp_mult_155(376);
partial_product_11(377) <= temp_mult_155(377);
partial_product_11(378) <= temp_mult_155(378);
partial_product_11(379) <= temp_mult_155(379);
partial_product_11(380) <= temp_mult_155(380);
partial_product_11(381) <= temp_mult_155(381);
partial_product_11(382) <= temp_mult_155(382);
partial_product_11(383) <= temp_mult_155(383);
partial_product_11(384) <= temp_mult_155(384);
partial_product_11(385) <= temp_mult_155(385);
partial_product_11(386) <= temp_mult_155(386);
partial_product_11(387) <= temp_mult_155(387);
partial_product_11(388) <= temp_mult_155(388);
partial_product_11(389) <= temp_mult_155(389);
partial_product_11(390) <= temp_mult_155(390);
partial_product_11(391) <= temp_mult_155(391);
partial_product_11(392) <= temp_mult_155(392);
partial_product_11(393) <= temp_mult_155(393);
partial_product_11(394) <= temp_mult_155(394);
partial_product_11(395) <= temp_mult_155(395);
partial_product_11(396) <= temp_mult_155(396);
partial_product_11(397) <= temp_mult_155(397);
partial_product_11(398) <= temp_mult_155(398);
partial_product_11(399) <= temp_mult_155(399);
partial_product_11(400) <= temp_mult_155(400);
partial_product_11(401) <= temp_mult_155(401);
partial_product_11(402) <= temp_mult_155(402);
partial_product_11(403) <= temp_mult_155(403);
partial_product_11(404) <= temp_mult_155(404);
partial_product_11(405) <= temp_mult_155(405);
partial_product_11(406) <= temp_mult_155(406);
partial_product_11(407) <= temp_mult_155(407);
partial_product_11(408) <= temp_mult_155(408);
partial_product_11(409) <= temp_mult_155(409);
partial_product_11(410) <= temp_mult_155(410);
partial_product_11(411) <= temp_mult_155(411);
partial_product_11(412) <= temp_mult_155(412);
partial_product_11(413) <= temp_mult_155(413);
partial_product_11(414) <= temp_mult_155(414);
partial_product_11(415) <= temp_mult_155(415);
partial_product_11(416) <= '0';
partial_product_11(417) <= '0';
partial_product_11(418) <= '0';
partial_product_11(419) <= '0';
partial_product_11(420) <= '0';
partial_product_11(421) <= '0';
partial_product_11(422) <= '0';
partial_product_11(423) <= '0';
partial_product_11(424) <= '0';
partial_product_11(425) <= '0';
partial_product_11(426) <= '0';
partial_product_11(427) <= '0';
partial_product_11(428) <= '0';
partial_product_11(429) <= '0';
partial_product_11(430) <= '0';
partial_product_11(431) <= '0';
partial_product_11(432) <= '0';
partial_product_11(433) <= '0';
partial_product_11(434) <= '0';
partial_product_11(435) <= '0';
partial_product_11(436) <= '0';
partial_product_11(437) <= '0';
partial_product_11(438) <= '0';
partial_product_11(439) <= '0';
partial_product_11(440) <= '0';
partial_product_11(441) <= '0';
partial_product_11(442) <= '0';
partial_product_11(443) <= '0';
partial_product_11(444) <= '0';
partial_product_11(445) <= '0';
partial_product_11(446) <= '0';
partial_product_11(447) <= '0';
partial_product_11(448) <= '0';
partial_product_11(449) <= '0';
partial_product_11(450) <= '0';
partial_product_11(451) <= '0';
partial_product_11(452) <= '0';
partial_product_11(453) <= '0';
partial_product_11(454) <= '0';
partial_product_11(455) <= '0';
partial_product_11(456) <= '0';
partial_product_11(457) <= '0';
partial_product_11(458) <= '0';
partial_product_11(459) <= '0';
partial_product_11(460) <= '0';
partial_product_11(461) <= '0';
partial_product_11(462) <= '0';
partial_product_11(463) <= '0';
partial_product_11(464) <= '0';
partial_product_11(465) <= '0';
partial_product_11(466) <= '0';
partial_product_11(467) <= '0';
partial_product_11(468) <= '0';
partial_product_11(469) <= '0';
partial_product_11(470) <= '0';
partial_product_11(471) <= '0';
partial_product_11(472) <= '0';
partial_product_11(473) <= '0';
partial_product_11(474) <= '0';
partial_product_11(475) <= '0';
partial_product_11(476) <= '0';
partial_product_11(477) <= '0';
partial_product_11(478) <= '0';
partial_product_11(479) <= '0';
partial_product_11(480) <= '0';
partial_product_11(481) <= '0';
partial_product_11(482) <= '0';
partial_product_11(483) <= '0';
partial_product_11(484) <= '0';
partial_product_11(485) <= '0';
partial_product_11(486) <= '0';
partial_product_11(487) <= '0';
partial_product_11(488) <= '0';
partial_product_11(489) <= '0';
partial_product_11(490) <= '0';
partial_product_11(491) <= '0';
partial_product_11(492) <= '0';
partial_product_11(493) <= '0';
partial_product_11(494) <= '0';
partial_product_11(495) <= '0';
partial_product_11(496) <= '0';
partial_product_11(497) <= '0';
partial_product_11(498) <= '0';
partial_product_11(499) <= '0';
partial_product_11(500) <= '0';
partial_product_11(501) <= '0';
partial_product_11(502) <= '0';
partial_product_11(503) <= '0';
partial_product_11(504) <= '0';
partial_product_11(505) <= '0';
partial_product_11(506) <= '0';
partial_product_11(507) <= '0';
partial_product_11(508) <= '0';
partial_product_11(509) <= '0';
partial_product_11(510) <= '0';
partial_product_11(511) <= '0';
partial_product_11(512) <= '0';
partial_product_12(0) <= '0';
partial_product_12(1) <= '0';
partial_product_12(2) <= '0';
partial_product_12(3) <= '0';
partial_product_12(4) <= '0';
partial_product_12(5) <= '0';
partial_product_12(6) <= '0';
partial_product_12(7) <= '0';
partial_product_12(8) <= '0';
partial_product_12(9) <= '0';
partial_product_12(10) <= '0';
partial_product_12(11) <= '0';
partial_product_12(12) <= '0';
partial_product_12(13) <= '0';
partial_product_12(14) <= '0';
partial_product_12(15) <= '0';
partial_product_12(16) <= '0';
partial_product_12(17) <= '0';
partial_product_12(18) <= '0';
partial_product_12(19) <= '0';
partial_product_12(20) <= '0';
partial_product_12(21) <= '0';
partial_product_12(22) <= '0';
partial_product_12(23) <= '0';
partial_product_12(24) <= '0';
partial_product_12(25) <= '0';
partial_product_12(26) <= '0';
partial_product_12(27) <= '0';
partial_product_12(28) <= '0';
partial_product_12(29) <= '0';
partial_product_12(30) <= '0';
partial_product_12(31) <= '0';
partial_product_12(32) <= '0';
partial_product_12(33) <= '0';
partial_product_12(34) <= '0';
partial_product_12(35) <= '0';
partial_product_12(36) <= '0';
partial_product_12(37) <= '0';
partial_product_12(38) <= '0';
partial_product_12(39) <= '0';
partial_product_12(40) <= '0';
partial_product_12(41) <= '0';
partial_product_12(42) <= '0';
partial_product_12(43) <= '0';
partial_product_12(44) <= '0';
partial_product_12(45) <= '0';
partial_product_12(46) <= '0';
partial_product_12(47) <= '0';
partial_product_12(48) <= '0';
partial_product_12(49) <= '0';
partial_product_12(50) <= '0';
partial_product_12(51) <= '0';
partial_product_12(52) <= '0';
partial_product_12(53) <= '0';
partial_product_12(54) <= '0';
partial_product_12(55) <= '0';
partial_product_12(56) <= '0';
partial_product_12(57) <= '0';
partial_product_12(58) <= '0';
partial_product_12(59) <= '0';
partial_product_12(60) <= '0';
partial_product_12(61) <= '0';
partial_product_12(62) <= '0';
partial_product_12(63) <= '0';
partial_product_12(64) <= '0';
partial_product_12(65) <= '0';
partial_product_12(66) <= '0';
partial_product_12(67) <= '0';
partial_product_12(68) <= '0';
partial_product_12(69) <= '0';
partial_product_12(70) <= '0';
partial_product_12(71) <= '0';
partial_product_12(72) <= '0';
partial_product_12(73) <= '0';
partial_product_12(74) <= '0';
partial_product_12(75) <= '0';
partial_product_12(76) <= '0';
partial_product_12(77) <= '0';
partial_product_12(78) <= '0';
partial_product_12(79) <= '0';
partial_product_12(80) <= '0';
partial_product_12(81) <= '0';
partial_product_12(82) <= '0';
partial_product_12(83) <= '0';
partial_product_12(84) <= '0';
partial_product_12(85) <= '0';
partial_product_12(86) <= '0';
partial_product_12(87) <= '0';
partial_product_12(88) <= '0';
partial_product_12(89) <= '0';
partial_product_12(90) <= '0';
partial_product_12(91) <= '0';
partial_product_12(92) <= '0';
partial_product_12(93) <= '0';
partial_product_12(94) <= '0';
partial_product_12(95) <= '0';
partial_product_12(96) <= '0';
partial_product_12(97) <= '0';
partial_product_12(98) <= '0';
partial_product_12(99) <= '0';
partial_product_12(100) <= '0';
partial_product_12(101) <= '0';
partial_product_12(102) <= '0';
partial_product_12(103) <= '0';
partial_product_12(104) <= '0';
partial_product_12(105) <= '0';
partial_product_12(106) <= '0';
partial_product_12(107) <= '0';
partial_product_12(108) <= '0';
partial_product_12(109) <= '0';
partial_product_12(110) <= '0';
partial_product_12(111) <= '0';
partial_product_12(112) <= '0';
partial_product_12(113) <= '0';
partial_product_12(114) <= '0';
partial_product_12(115) <= '0';
partial_product_12(116) <= '0';
partial_product_12(117) <= '0';
partial_product_12(118) <= '0';
partial_product_12(119) <= '0';
partial_product_12(120) <= temp_mult_40(120);
partial_product_12(121) <= temp_mult_40(121);
partial_product_12(122) <= temp_mult_40(122);
partial_product_12(123) <= temp_mult_40(123);
partial_product_12(124) <= temp_mult_40(124);
partial_product_12(125) <= temp_mult_40(125);
partial_product_12(126) <= temp_mult_40(126);
partial_product_12(127) <= temp_mult_40(127);
partial_product_12(128) <= temp_mult_40(128);
partial_product_12(129) <= temp_mult_40(129);
partial_product_12(130) <= temp_mult_40(130);
partial_product_12(131) <= temp_mult_40(131);
partial_product_12(132) <= temp_mult_40(132);
partial_product_12(133) <= temp_mult_40(133);
partial_product_12(134) <= temp_mult_40(134);
partial_product_12(135) <= temp_mult_40(135);
partial_product_12(136) <= temp_mult_40(136);
partial_product_12(137) <= temp_mult_40(137);
partial_product_12(138) <= temp_mult_40(138);
partial_product_12(139) <= temp_mult_40(139);
partial_product_12(140) <= temp_mult_40(140);
partial_product_12(141) <= temp_mult_40(141);
partial_product_12(142) <= temp_mult_40(142);
partial_product_12(143) <= temp_mult_40(143);
partial_product_12(144) <= temp_mult_40(144);
partial_product_12(145) <= temp_mult_40(145);
partial_product_12(146) <= temp_mult_40(146);
partial_product_12(147) <= temp_mult_40(147);
partial_product_12(148) <= temp_mult_40(148);
partial_product_12(149) <= temp_mult_40(149);
partial_product_12(150) <= temp_mult_40(150);
partial_product_12(151) <= temp_mult_40(151);
partial_product_12(152) <= temp_mult_40(152);
partial_product_12(153) <= temp_mult_40(153);
partial_product_12(154) <= temp_mult_40(154);
partial_product_12(155) <= temp_mult_40(155);
partial_product_12(156) <= temp_mult_40(156);
partial_product_12(157) <= temp_mult_40(157);
partial_product_12(158) <= temp_mult_40(158);
partial_product_12(159) <= temp_mult_40(159);
partial_product_12(160) <= temp_mult_40(160);
partial_product_12(161) <= temp_mult_49(161);
partial_product_12(162) <= temp_mult_49(162);
partial_product_12(163) <= temp_mult_49(163);
partial_product_12(164) <= temp_mult_49(164);
partial_product_12(165) <= temp_mult_49(165);
partial_product_12(166) <= temp_mult_49(166);
partial_product_12(167) <= temp_mult_49(167);
partial_product_12(168) <= temp_mult_49(168);
partial_product_12(169) <= temp_mult_49(169);
partial_product_12(170) <= temp_mult_49(170);
partial_product_12(171) <= temp_mult_49(171);
partial_product_12(172) <= temp_mult_49(172);
partial_product_12(173) <= temp_mult_49(173);
partial_product_12(174) <= temp_mult_49(174);
partial_product_12(175) <= temp_mult_49(175);
partial_product_12(176) <= temp_mult_49(176);
partial_product_12(177) <= temp_mult_49(177);
partial_product_12(178) <= temp_mult_49(178);
partial_product_12(179) <= temp_mult_49(179);
partial_product_12(180) <= temp_mult_49(180);
partial_product_12(181) <= temp_mult_49(181);
partial_product_12(182) <= temp_mult_49(182);
partial_product_12(183) <= temp_mult_49(183);
partial_product_12(184) <= temp_mult_49(184);
partial_product_12(185) <= temp_mult_49(185);
partial_product_12(186) <= temp_mult_49(186);
partial_product_12(187) <= temp_mult_49(187);
partial_product_12(188) <= temp_mult_49(188);
partial_product_12(189) <= temp_mult_49(189);
partial_product_12(190) <= temp_mult_49(190);
partial_product_12(191) <= temp_mult_49(191);
partial_product_12(192) <= temp_mult_49(192);
partial_product_12(193) <= temp_mult_49(193);
partial_product_12(194) <= temp_mult_49(194);
partial_product_12(195) <= temp_mult_49(195);
partial_product_12(196) <= temp_mult_49(196);
partial_product_12(197) <= temp_mult_49(197);
partial_product_12(198) <= temp_mult_49(198);
partial_product_12(199) <= temp_mult_49(199);
partial_product_12(200) <= temp_mult_49(200);
partial_product_12(201) <= temp_mult_49(201);
partial_product_12(202) <= temp_mult_58(202);
partial_product_12(203) <= temp_mult_58(203);
partial_product_12(204) <= temp_mult_58(204);
partial_product_12(205) <= temp_mult_58(205);
partial_product_12(206) <= temp_mult_58(206);
partial_product_12(207) <= temp_mult_58(207);
partial_product_12(208) <= temp_mult_58(208);
partial_product_12(209) <= temp_mult_58(209);
partial_product_12(210) <= temp_mult_58(210);
partial_product_12(211) <= temp_mult_58(211);
partial_product_12(212) <= temp_mult_58(212);
partial_product_12(213) <= temp_mult_58(213);
partial_product_12(214) <= temp_mult_58(214);
partial_product_12(215) <= temp_mult_58(215);
partial_product_12(216) <= temp_mult_58(216);
partial_product_12(217) <= temp_mult_58(217);
partial_product_12(218) <= temp_mult_58(218);
partial_product_12(219) <= temp_mult_58(219);
partial_product_12(220) <= temp_mult_58(220);
partial_product_12(221) <= temp_mult_58(221);
partial_product_12(222) <= temp_mult_58(222);
partial_product_12(223) <= temp_mult_58(223);
partial_product_12(224) <= temp_mult_58(224);
partial_product_12(225) <= temp_mult_58(225);
partial_product_12(226) <= temp_mult_58(226);
partial_product_12(227) <= temp_mult_58(227);
partial_product_12(228) <= temp_mult_58(228);
partial_product_12(229) <= temp_mult_58(229);
partial_product_12(230) <= temp_mult_58(230);
partial_product_12(231) <= temp_mult_58(231);
partial_product_12(232) <= temp_mult_58(232);
partial_product_12(233) <= temp_mult_58(233);
partial_product_12(234) <= temp_mult_58(234);
partial_product_12(235) <= temp_mult_58(235);
partial_product_12(236) <= temp_mult_58(236);
partial_product_12(237) <= temp_mult_58(237);
partial_product_12(238) <= temp_mult_58(238);
partial_product_12(239) <= temp_mult_58(239);
partial_product_12(240) <= temp_mult_58(240);
partial_product_12(241) <= temp_mult_58(241);
partial_product_12(242) <= temp_mult_58(242);
partial_product_12(243) <= temp_mult_67(243);
partial_product_12(244) <= temp_mult_67(244);
partial_product_12(245) <= temp_mult_67(245);
partial_product_12(246) <= temp_mult_67(246);
partial_product_12(247) <= temp_mult_67(247);
partial_product_12(248) <= temp_mult_67(248);
partial_product_12(249) <= temp_mult_67(249);
partial_product_12(250) <= temp_mult_67(250);
partial_product_12(251) <= temp_mult_67(251);
partial_product_12(252) <= temp_mult_67(252);
partial_product_12(253) <= temp_mult_67(253);
partial_product_12(254) <= temp_mult_67(254);
partial_product_12(255) <= temp_mult_67(255);
partial_product_12(256) <= temp_mult_67(256);
partial_product_12(257) <= temp_mult_67(257);
partial_product_12(258) <= temp_mult_67(258);
partial_product_12(259) <= temp_mult_67(259);
partial_product_12(260) <= temp_mult_67(260);
partial_product_12(261) <= temp_mult_67(261);
partial_product_12(262) <= temp_mult_67(262);
partial_product_12(263) <= temp_mult_67(263);
partial_product_12(264) <= temp_mult_67(264);
partial_product_12(265) <= temp_mult_67(265);
partial_product_12(266) <= temp_mult_67(266);
partial_product_12(267) <= temp_mult_67(267);
partial_product_12(268) <= temp_mult_67(268);
partial_product_12(269) <= temp_mult_67(269);
partial_product_12(270) <= temp_mult_67(270);
partial_product_12(271) <= temp_mult_67(271);
partial_product_12(272) <= temp_mult_67(272);
partial_product_12(273) <= temp_mult_67(273);
partial_product_12(274) <= temp_mult_67(274);
partial_product_12(275) <= temp_mult_67(275);
partial_product_12(276) <= temp_mult_67(276);
partial_product_12(277) <= temp_mult_67(277);
partial_product_12(278) <= temp_mult_67(278);
partial_product_12(279) <= temp_mult_67(279);
partial_product_12(280) <= temp_mult_67(280);
partial_product_12(281) <= temp_mult_67(281);
partial_product_12(282) <= temp_mult_67(282);
partial_product_12(283) <= temp_mult_67(283);
partial_product_12(284) <= temp_mult_76(284);
partial_product_12(285) <= temp_mult_76(285);
partial_product_12(286) <= temp_mult_76(286);
partial_product_12(287) <= temp_mult_76(287);
partial_product_12(288) <= temp_mult_76(288);
partial_product_12(289) <= temp_mult_76(289);
partial_product_12(290) <= temp_mult_76(290);
partial_product_12(291) <= temp_mult_76(291);
partial_product_12(292) <= temp_mult_76(292);
partial_product_12(293) <= temp_mult_76(293);
partial_product_12(294) <= temp_mult_76(294);
partial_product_12(295) <= temp_mult_76(295);
partial_product_12(296) <= temp_mult_76(296);
partial_product_12(297) <= temp_mult_76(297);
partial_product_12(298) <= temp_mult_76(298);
partial_product_12(299) <= temp_mult_76(299);
partial_product_12(300) <= temp_mult_76(300);
partial_product_12(301) <= temp_mult_76(301);
partial_product_12(302) <= temp_mult_76(302);
partial_product_12(303) <= temp_mult_76(303);
partial_product_12(304) <= temp_mult_76(304);
partial_product_12(305) <= temp_mult_76(305);
partial_product_12(306) <= temp_mult_76(306);
partial_product_12(307) <= temp_mult_76(307);
partial_product_12(308) <= temp_mult_76(308);
partial_product_12(309) <= temp_mult_76(309);
partial_product_12(310) <= temp_mult_76(310);
partial_product_12(311) <= temp_mult_76(311);
partial_product_12(312) <= temp_mult_76(312);
partial_product_12(313) <= temp_mult_76(313);
partial_product_12(314) <= temp_mult_76(314);
partial_product_12(315) <= temp_mult_76(315);
partial_product_12(316) <= temp_mult_76(316);
partial_product_12(317) <= temp_mult_76(317);
partial_product_12(318) <= temp_mult_76(318);
partial_product_12(319) <= temp_mult_76(319);
partial_product_12(320) <= temp_mult_76(320);
partial_product_12(321) <= temp_mult_76(321);
partial_product_12(322) <= temp_mult_76(322);
partial_product_12(323) <= temp_mult_76(323);
partial_product_12(324) <= temp_mult_76(324);
partial_product_12(325) <= '0';
partial_product_12(326) <= '0';
partial_product_12(327) <= temp_mult_111(327);
partial_product_12(328) <= temp_mult_111(328);
partial_product_12(329) <= temp_mult_111(329);
partial_product_12(330) <= temp_mult_111(330);
partial_product_12(331) <= temp_mult_111(331);
partial_product_12(332) <= temp_mult_111(332);
partial_product_12(333) <= temp_mult_111(333);
partial_product_12(334) <= temp_mult_111(334);
partial_product_12(335) <= temp_mult_111(335);
partial_product_12(336) <= temp_mult_111(336);
partial_product_12(337) <= temp_mult_111(337);
partial_product_12(338) <= temp_mult_111(338);
partial_product_12(339) <= temp_mult_111(339);
partial_product_12(340) <= temp_mult_111(340);
partial_product_12(341) <= temp_mult_111(341);
partial_product_12(342) <= temp_mult_111(342);
partial_product_12(343) <= temp_mult_111(343);
partial_product_12(344) <= temp_mult_111(344);
partial_product_12(345) <= temp_mult_111(345);
partial_product_12(346) <= temp_mult_111(346);
partial_product_12(347) <= temp_mult_111(347);
partial_product_12(348) <= temp_mult_111(348);
partial_product_12(349) <= temp_mult_111(349);
partial_product_12(350) <= temp_mult_111(350);
partial_product_12(351) <= temp_mult_111(351);
partial_product_12(352) <= temp_mult_111(352);
partial_product_12(353) <= temp_mult_111(353);
partial_product_12(354) <= temp_mult_111(354);
partial_product_12(355) <= temp_mult_111(355);
partial_product_12(356) <= temp_mult_111(356);
partial_product_12(357) <= temp_mult_111(357);
partial_product_12(358) <= temp_mult_111(358);
partial_product_12(359) <= temp_mult_111(359);
partial_product_12(360) <= temp_mult_111(360);
partial_product_12(361) <= temp_mult_111(361);
partial_product_12(362) <= temp_mult_111(362);
partial_product_12(363) <= temp_mult_111(363);
partial_product_12(364) <= temp_mult_111(364);
partial_product_12(365) <= temp_mult_111(365);
partial_product_12(366) <= temp_mult_111(366);
partial_product_12(367) <= temp_mult_111(367);
partial_product_12(368) <= '0';
partial_product_12(369) <= '0';
partial_product_12(370) <= '0';
partial_product_12(371) <= '0';
partial_product_12(372) <= '0';
partial_product_12(373) <= '0';
partial_product_12(374) <= '0';
partial_product_12(375) <= '0';
partial_product_12(376) <= '0';
partial_product_12(377) <= '0';
partial_product_12(378) <= '0';
partial_product_12(379) <= '0';
partial_product_12(380) <= '0';
partial_product_12(381) <= '0';
partial_product_12(382) <= '0';
partial_product_12(383) <= '0';
partial_product_12(384) <= '0';
partial_product_12(385) <= '0';
partial_product_12(386) <= '0';
partial_product_12(387) <= '0';
partial_product_12(388) <= '0';
partial_product_12(389) <= '0';
partial_product_12(390) <= '0';
partial_product_12(391) <= '0';
partial_product_12(392) <= '0';
partial_product_12(393) <= '0';
partial_product_12(394) <= '0';
partial_product_12(395) <= '0';
partial_product_12(396) <= '0';
partial_product_12(397) <= '0';
partial_product_12(398) <= '0';
partial_product_12(399) <= '0';
partial_product_12(400) <= '0';
partial_product_12(401) <= '0';
partial_product_12(402) <= '0';
partial_product_12(403) <= '0';
partial_product_12(404) <= '0';
partial_product_12(405) <= '0';
partial_product_12(406) <= '0';
partial_product_12(407) <= '0';
partial_product_12(408) <= '0';
partial_product_12(409) <= '0';
partial_product_12(410) <= '0';
partial_product_12(411) <= '0';
partial_product_12(412) <= '0';
partial_product_12(413) <= '0';
partial_product_12(414) <= '0';
partial_product_12(415) <= '0';
partial_product_12(416) <= '0';
partial_product_12(417) <= '0';
partial_product_12(418) <= '0';
partial_product_12(419) <= '0';
partial_product_12(420) <= '0';
partial_product_12(421) <= '0';
partial_product_12(422) <= '0';
partial_product_12(423) <= '0';
partial_product_12(424) <= '0';
partial_product_12(425) <= '0';
partial_product_12(426) <= '0';
partial_product_12(427) <= '0';
partial_product_12(428) <= '0';
partial_product_12(429) <= '0';
partial_product_12(430) <= '0';
partial_product_12(431) <= '0';
partial_product_12(432) <= '0';
partial_product_12(433) <= '0';
partial_product_12(434) <= '0';
partial_product_12(435) <= '0';
partial_product_12(436) <= '0';
partial_product_12(437) <= '0';
partial_product_12(438) <= '0';
partial_product_12(439) <= '0';
partial_product_12(440) <= '0';
partial_product_12(441) <= '0';
partial_product_12(442) <= '0';
partial_product_12(443) <= '0';
partial_product_12(444) <= '0';
partial_product_12(445) <= '0';
partial_product_12(446) <= '0';
partial_product_12(447) <= '0';
partial_product_12(448) <= '0';
partial_product_12(449) <= '0';
partial_product_12(450) <= '0';
partial_product_12(451) <= '0';
partial_product_12(452) <= '0';
partial_product_12(453) <= '0';
partial_product_12(454) <= '0';
partial_product_12(455) <= '0';
partial_product_12(456) <= '0';
partial_product_12(457) <= '0';
partial_product_12(458) <= '0';
partial_product_12(459) <= '0';
partial_product_12(460) <= '0';
partial_product_12(461) <= '0';
partial_product_12(462) <= '0';
partial_product_12(463) <= '0';
partial_product_12(464) <= '0';
partial_product_12(465) <= '0';
partial_product_12(466) <= '0';
partial_product_12(467) <= '0';
partial_product_12(468) <= '0';
partial_product_12(469) <= '0';
partial_product_12(470) <= '0';
partial_product_12(471) <= '0';
partial_product_12(472) <= '0';
partial_product_12(473) <= '0';
partial_product_12(474) <= '0';
partial_product_12(475) <= '0';
partial_product_12(476) <= '0';
partial_product_12(477) <= '0';
partial_product_12(478) <= '0';
partial_product_12(479) <= '0';
partial_product_12(480) <= '0';
partial_product_12(481) <= '0';
partial_product_12(482) <= '0';
partial_product_12(483) <= '0';
partial_product_12(484) <= '0';
partial_product_12(485) <= '0';
partial_product_12(486) <= '0';
partial_product_12(487) <= '0';
partial_product_12(488) <= '0';
partial_product_12(489) <= '0';
partial_product_12(490) <= '0';
partial_product_12(491) <= '0';
partial_product_12(492) <= '0';
partial_product_12(493) <= '0';
partial_product_12(494) <= '0';
partial_product_12(495) <= '0';
partial_product_12(496) <= '0';
partial_product_12(497) <= '0';
partial_product_12(498) <= '0';
partial_product_12(499) <= '0';
partial_product_12(500) <= '0';
partial_product_12(501) <= '0';
partial_product_12(502) <= '0';
partial_product_12(503) <= '0';
partial_product_12(504) <= '0';
partial_product_12(505) <= '0';
partial_product_12(506) <= '0';
partial_product_12(507) <= '0';
partial_product_12(508) <= '0';
partial_product_12(509) <= '0';
partial_product_12(510) <= '0';
partial_product_12(511) <= '0';
partial_product_12(512) <= '0';
partial_product_13(0) <= '0';
partial_product_13(1) <= '0';
partial_product_13(2) <= '0';
partial_product_13(3) <= '0';
partial_product_13(4) <= '0';
partial_product_13(5) <= '0';
partial_product_13(6) <= '0';
partial_product_13(7) <= '0';
partial_product_13(8) <= '0';
partial_product_13(9) <= '0';
partial_product_13(10) <= '0';
partial_product_13(11) <= '0';
partial_product_13(12) <= '0';
partial_product_13(13) <= '0';
partial_product_13(14) <= '0';
partial_product_13(15) <= '0';
partial_product_13(16) <= '0';
partial_product_13(17) <= '0';
partial_product_13(18) <= '0';
partial_product_13(19) <= '0';
partial_product_13(20) <= '0';
partial_product_13(21) <= '0';
partial_product_13(22) <= '0';
partial_product_13(23) <= '0';
partial_product_13(24) <= '0';
partial_product_13(25) <= '0';
partial_product_13(26) <= '0';
partial_product_13(27) <= '0';
partial_product_13(28) <= '0';
partial_product_13(29) <= '0';
partial_product_13(30) <= '0';
partial_product_13(31) <= '0';
partial_product_13(32) <= '0';
partial_product_13(33) <= '0';
partial_product_13(34) <= '0';
partial_product_13(35) <= '0';
partial_product_13(36) <= '0';
partial_product_13(37) <= '0';
partial_product_13(38) <= '0';
partial_product_13(39) <= '0';
partial_product_13(40) <= '0';
partial_product_13(41) <= '0';
partial_product_13(42) <= '0';
partial_product_13(43) <= '0';
partial_product_13(44) <= '0';
partial_product_13(45) <= '0';
partial_product_13(46) <= '0';
partial_product_13(47) <= '0';
partial_product_13(48) <= '0';
partial_product_13(49) <= '0';
partial_product_13(50) <= '0';
partial_product_13(51) <= '0';
partial_product_13(52) <= '0';
partial_product_13(53) <= '0';
partial_product_13(54) <= '0';
partial_product_13(55) <= '0';
partial_product_13(56) <= '0';
partial_product_13(57) <= '0';
partial_product_13(58) <= '0';
partial_product_13(59) <= '0';
partial_product_13(60) <= '0';
partial_product_13(61) <= '0';
partial_product_13(62) <= '0';
partial_product_13(63) <= '0';
partial_product_13(64) <= '0';
partial_product_13(65) <= '0';
partial_product_13(66) <= '0';
partial_product_13(67) <= '0';
partial_product_13(68) <= '0';
partial_product_13(69) <= '0';
partial_product_13(70) <= '0';
partial_product_13(71) <= '0';
partial_product_13(72) <= '0';
partial_product_13(73) <= '0';
partial_product_13(74) <= '0';
partial_product_13(75) <= '0';
partial_product_13(76) <= '0';
partial_product_13(77) <= '0';
partial_product_13(78) <= '0';
partial_product_13(79) <= '0';
partial_product_13(80) <= '0';
partial_product_13(81) <= '0';
partial_product_13(82) <= '0';
partial_product_13(83) <= '0';
partial_product_13(84) <= '0';
partial_product_13(85) <= '0';
partial_product_13(86) <= '0';
partial_product_13(87) <= '0';
partial_product_13(88) <= '0';
partial_product_13(89) <= '0';
partial_product_13(90) <= '0';
partial_product_13(91) <= '0';
partial_product_13(92) <= '0';
partial_product_13(93) <= '0';
partial_product_13(94) <= '0';
partial_product_13(95) <= '0';
partial_product_13(96) <= '0';
partial_product_13(97) <= '0';
partial_product_13(98) <= '0';
partial_product_13(99) <= '0';
partial_product_13(100) <= '0';
partial_product_13(101) <= '0';
partial_product_13(102) <= '0';
partial_product_13(103) <= '0';
partial_product_13(104) <= '0';
partial_product_13(105) <= '0';
partial_product_13(106) <= '0';
partial_product_13(107) <= '0';
partial_product_13(108) <= '0';
partial_product_13(109) <= '0';
partial_product_13(110) <= '0';
partial_product_13(111) <= '0';
partial_product_13(112) <= '0';
partial_product_13(113) <= '0';
partial_product_13(114) <= '0';
partial_product_13(115) <= '0';
partial_product_13(116) <= '0';
partial_product_13(117) <= '0';
partial_product_13(118) <= '0';
partial_product_13(119) <= '0';
partial_product_13(120) <= '0';
partial_product_13(121) <= '0';
partial_product_13(122) <= '0';
partial_product_13(123) <= '0';
partial_product_13(124) <= '0';
partial_product_13(125) <= '0';
partial_product_13(126) <= '0';
partial_product_13(127) <= '0';
partial_product_13(128) <= '0';
partial_product_13(129) <= '0';
partial_product_13(130) <= '0';
partial_product_13(131) <= '0';
partial_product_13(132) <= '0';
partial_product_13(133) <= '0';
partial_product_13(134) <= '0';
partial_product_13(135) <= '0';
partial_product_13(136) <= temp_mult_80(136);
partial_product_13(137) <= temp_mult_80(137);
partial_product_13(138) <= temp_mult_80(138);
partial_product_13(139) <= temp_mult_80(139);
partial_product_13(140) <= temp_mult_80(140);
partial_product_13(141) <= temp_mult_80(141);
partial_product_13(142) <= temp_mult_80(142);
partial_product_13(143) <= temp_mult_80(143);
partial_product_13(144) <= temp_mult_80(144);
partial_product_13(145) <= temp_mult_80(145);
partial_product_13(146) <= temp_mult_80(146);
partial_product_13(147) <= temp_mult_80(147);
partial_product_13(148) <= temp_mult_80(148);
partial_product_13(149) <= temp_mult_80(149);
partial_product_13(150) <= temp_mult_80(150);
partial_product_13(151) <= temp_mult_80(151);
partial_product_13(152) <= temp_mult_80(152);
partial_product_13(153) <= temp_mult_80(153);
partial_product_13(154) <= temp_mult_80(154);
partial_product_13(155) <= temp_mult_80(155);
partial_product_13(156) <= temp_mult_80(156);
partial_product_13(157) <= temp_mult_80(157);
partial_product_13(158) <= temp_mult_80(158);
partial_product_13(159) <= temp_mult_80(159);
partial_product_13(160) <= temp_mult_80(160);
partial_product_13(161) <= temp_mult_80(161);
partial_product_13(162) <= temp_mult_80(162);
partial_product_13(163) <= temp_mult_80(163);
partial_product_13(164) <= temp_mult_80(164);
partial_product_13(165) <= temp_mult_80(165);
partial_product_13(166) <= temp_mult_80(166);
partial_product_13(167) <= temp_mult_80(167);
partial_product_13(168) <= temp_mult_80(168);
partial_product_13(169) <= temp_mult_80(169);
partial_product_13(170) <= temp_mult_80(170);
partial_product_13(171) <= temp_mult_80(171);
partial_product_13(172) <= temp_mult_80(172);
partial_product_13(173) <= temp_mult_80(173);
partial_product_13(174) <= temp_mult_80(174);
partial_product_13(175) <= temp_mult_80(175);
partial_product_13(176) <= temp_mult_80(176);
partial_product_13(177) <= temp_mult_89(177);
partial_product_13(178) <= temp_mult_89(178);
partial_product_13(179) <= temp_mult_89(179);
partial_product_13(180) <= temp_mult_89(180);
partial_product_13(181) <= temp_mult_89(181);
partial_product_13(182) <= temp_mult_89(182);
partial_product_13(183) <= temp_mult_89(183);
partial_product_13(184) <= temp_mult_89(184);
partial_product_13(185) <= temp_mult_89(185);
partial_product_13(186) <= temp_mult_89(186);
partial_product_13(187) <= temp_mult_89(187);
partial_product_13(188) <= temp_mult_89(188);
partial_product_13(189) <= temp_mult_89(189);
partial_product_13(190) <= temp_mult_89(190);
partial_product_13(191) <= temp_mult_89(191);
partial_product_13(192) <= temp_mult_89(192);
partial_product_13(193) <= temp_mult_89(193);
partial_product_13(194) <= temp_mult_89(194);
partial_product_13(195) <= temp_mult_89(195);
partial_product_13(196) <= temp_mult_89(196);
partial_product_13(197) <= temp_mult_89(197);
partial_product_13(198) <= temp_mult_89(198);
partial_product_13(199) <= temp_mult_89(199);
partial_product_13(200) <= temp_mult_89(200);
partial_product_13(201) <= temp_mult_89(201);
partial_product_13(202) <= temp_mult_89(202);
partial_product_13(203) <= temp_mult_89(203);
partial_product_13(204) <= temp_mult_89(204);
partial_product_13(205) <= temp_mult_89(205);
partial_product_13(206) <= temp_mult_89(206);
partial_product_13(207) <= temp_mult_89(207);
partial_product_13(208) <= temp_mult_89(208);
partial_product_13(209) <= temp_mult_89(209);
partial_product_13(210) <= temp_mult_89(210);
partial_product_13(211) <= temp_mult_89(211);
partial_product_13(212) <= temp_mult_89(212);
partial_product_13(213) <= temp_mult_89(213);
partial_product_13(214) <= temp_mult_89(214);
partial_product_13(215) <= temp_mult_89(215);
partial_product_13(216) <= temp_mult_89(216);
partial_product_13(217) <= temp_mult_89(217);
partial_product_13(218) <= temp_mult_98(218);
partial_product_13(219) <= temp_mult_98(219);
partial_product_13(220) <= temp_mult_98(220);
partial_product_13(221) <= temp_mult_98(221);
partial_product_13(222) <= temp_mult_98(222);
partial_product_13(223) <= temp_mult_98(223);
partial_product_13(224) <= temp_mult_98(224);
partial_product_13(225) <= temp_mult_98(225);
partial_product_13(226) <= temp_mult_98(226);
partial_product_13(227) <= temp_mult_98(227);
partial_product_13(228) <= temp_mult_98(228);
partial_product_13(229) <= temp_mult_98(229);
partial_product_13(230) <= temp_mult_98(230);
partial_product_13(231) <= temp_mult_98(231);
partial_product_13(232) <= temp_mult_98(232);
partial_product_13(233) <= temp_mult_98(233);
partial_product_13(234) <= temp_mult_98(234);
partial_product_13(235) <= temp_mult_98(235);
partial_product_13(236) <= temp_mult_98(236);
partial_product_13(237) <= temp_mult_98(237);
partial_product_13(238) <= temp_mult_98(238);
partial_product_13(239) <= temp_mult_98(239);
partial_product_13(240) <= temp_mult_98(240);
partial_product_13(241) <= temp_mult_98(241);
partial_product_13(242) <= temp_mult_98(242);
partial_product_13(243) <= temp_mult_98(243);
partial_product_13(244) <= temp_mult_98(244);
partial_product_13(245) <= temp_mult_98(245);
partial_product_13(246) <= temp_mult_98(246);
partial_product_13(247) <= temp_mult_98(247);
partial_product_13(248) <= temp_mult_98(248);
partial_product_13(249) <= temp_mult_98(249);
partial_product_13(250) <= temp_mult_98(250);
partial_product_13(251) <= temp_mult_98(251);
partial_product_13(252) <= temp_mult_98(252);
partial_product_13(253) <= temp_mult_98(253);
partial_product_13(254) <= temp_mult_98(254);
partial_product_13(255) <= temp_mult_98(255);
partial_product_13(256) <= temp_mult_98(256);
partial_product_13(257) <= temp_mult_98(257);
partial_product_13(258) <= temp_mult_98(258);
partial_product_13(259) <= temp_mult_107(259);
partial_product_13(260) <= temp_mult_107(260);
partial_product_13(261) <= temp_mult_107(261);
partial_product_13(262) <= temp_mult_107(262);
partial_product_13(263) <= temp_mult_107(263);
partial_product_13(264) <= temp_mult_107(264);
partial_product_13(265) <= temp_mult_107(265);
partial_product_13(266) <= temp_mult_107(266);
partial_product_13(267) <= temp_mult_107(267);
partial_product_13(268) <= temp_mult_107(268);
partial_product_13(269) <= temp_mult_107(269);
partial_product_13(270) <= temp_mult_107(270);
partial_product_13(271) <= temp_mult_107(271);
partial_product_13(272) <= temp_mult_107(272);
partial_product_13(273) <= temp_mult_107(273);
partial_product_13(274) <= temp_mult_107(274);
partial_product_13(275) <= temp_mult_107(275);
partial_product_13(276) <= temp_mult_107(276);
partial_product_13(277) <= temp_mult_107(277);
partial_product_13(278) <= temp_mult_107(278);
partial_product_13(279) <= temp_mult_107(279);
partial_product_13(280) <= temp_mult_107(280);
partial_product_13(281) <= temp_mult_107(281);
partial_product_13(282) <= temp_mult_107(282);
partial_product_13(283) <= temp_mult_107(283);
partial_product_13(284) <= temp_mult_107(284);
partial_product_13(285) <= temp_mult_107(285);
partial_product_13(286) <= temp_mult_107(286);
partial_product_13(287) <= temp_mult_107(287);
partial_product_13(288) <= temp_mult_107(288);
partial_product_13(289) <= temp_mult_107(289);
partial_product_13(290) <= temp_mult_107(290);
partial_product_13(291) <= temp_mult_107(291);
partial_product_13(292) <= temp_mult_107(292);
partial_product_13(293) <= temp_mult_107(293);
partial_product_13(294) <= temp_mult_107(294);
partial_product_13(295) <= temp_mult_107(295);
partial_product_13(296) <= temp_mult_107(296);
partial_product_13(297) <= temp_mult_107(297);
partial_product_13(298) <= temp_mult_107(298);
partial_product_13(299) <= temp_mult_107(299);
partial_product_13(300) <= temp_mult_116(300);
partial_product_13(301) <= temp_mult_116(301);
partial_product_13(302) <= temp_mult_116(302);
partial_product_13(303) <= temp_mult_116(303);
partial_product_13(304) <= temp_mult_116(304);
partial_product_13(305) <= temp_mult_116(305);
partial_product_13(306) <= temp_mult_116(306);
partial_product_13(307) <= temp_mult_116(307);
partial_product_13(308) <= temp_mult_116(308);
partial_product_13(309) <= temp_mult_116(309);
partial_product_13(310) <= temp_mult_116(310);
partial_product_13(311) <= temp_mult_116(311);
partial_product_13(312) <= temp_mult_116(312);
partial_product_13(313) <= temp_mult_116(313);
partial_product_13(314) <= temp_mult_116(314);
partial_product_13(315) <= temp_mult_116(315);
partial_product_13(316) <= temp_mult_116(316);
partial_product_13(317) <= temp_mult_116(317);
partial_product_13(318) <= temp_mult_116(318);
partial_product_13(319) <= temp_mult_116(319);
partial_product_13(320) <= temp_mult_116(320);
partial_product_13(321) <= temp_mult_116(321);
partial_product_13(322) <= temp_mult_116(322);
partial_product_13(323) <= temp_mult_116(323);
partial_product_13(324) <= temp_mult_116(324);
partial_product_13(325) <= temp_mult_116(325);
partial_product_13(326) <= temp_mult_116(326);
partial_product_13(327) <= temp_mult_116(327);
partial_product_13(328) <= temp_mult_116(328);
partial_product_13(329) <= temp_mult_116(329);
partial_product_13(330) <= temp_mult_116(330);
partial_product_13(331) <= temp_mult_116(331);
partial_product_13(332) <= temp_mult_116(332);
partial_product_13(333) <= temp_mult_116(333);
partial_product_13(334) <= temp_mult_116(334);
partial_product_13(335) <= temp_mult_116(335);
partial_product_13(336) <= temp_mult_116(336);
partial_product_13(337) <= temp_mult_116(337);
partial_product_13(338) <= temp_mult_116(338);
partial_product_13(339) <= temp_mult_116(339);
partial_product_13(340) <= temp_mult_116(340);
partial_product_13(341) <= temp_mult_145(341);
partial_product_13(342) <= temp_mult_145(342);
partial_product_13(343) <= temp_mult_145(343);
partial_product_13(344) <= temp_mult_145(344);
partial_product_13(345) <= temp_mult_145(345);
partial_product_13(346) <= temp_mult_145(346);
partial_product_13(347) <= temp_mult_145(347);
partial_product_13(348) <= temp_mult_145(348);
partial_product_13(349) <= temp_mult_145(349);
partial_product_13(350) <= temp_mult_145(350);
partial_product_13(351) <= temp_mult_145(351);
partial_product_13(352) <= temp_mult_145(352);
partial_product_13(353) <= temp_mult_145(353);
partial_product_13(354) <= temp_mult_145(354);
partial_product_13(355) <= temp_mult_145(355);
partial_product_13(356) <= temp_mult_145(356);
partial_product_13(357) <= temp_mult_145(357);
partial_product_13(358) <= temp_mult_145(358);
partial_product_13(359) <= temp_mult_145(359);
partial_product_13(360) <= temp_mult_145(360);
partial_product_13(361) <= temp_mult_145(361);
partial_product_13(362) <= temp_mult_145(362);
partial_product_13(363) <= temp_mult_145(363);
partial_product_13(364) <= temp_mult_145(364);
partial_product_13(365) <= temp_mult_145(365);
partial_product_13(366) <= temp_mult_145(366);
partial_product_13(367) <= temp_mult_145(367);
partial_product_13(368) <= temp_mult_145(368);
partial_product_13(369) <= temp_mult_145(369);
partial_product_13(370) <= temp_mult_145(370);
partial_product_13(371) <= temp_mult_145(371);
partial_product_13(372) <= temp_mult_145(372);
partial_product_13(373) <= temp_mult_145(373);
partial_product_13(374) <= temp_mult_145(374);
partial_product_13(375) <= temp_mult_145(375);
partial_product_13(376) <= temp_mult_145(376);
partial_product_13(377) <= temp_mult_145(377);
partial_product_13(378) <= temp_mult_145(378);
partial_product_13(379) <= temp_mult_145(379);
partial_product_13(380) <= temp_mult_145(380);
partial_product_13(381) <= temp_mult_145(381);
partial_product_13(382) <= '0';
partial_product_13(383) <= '0';
partial_product_13(384) <= '0';
partial_product_13(385) <= '0';
partial_product_13(386) <= '0';
partial_product_13(387) <= '0';
partial_product_13(388) <= '0';
partial_product_13(389) <= '0';
partial_product_13(390) <= '0';
partial_product_13(391) <= '0';
partial_product_13(392) <= '0';
partial_product_13(393) <= '0';
partial_product_13(394) <= '0';
partial_product_13(395) <= '0';
partial_product_13(396) <= '0';
partial_product_13(397) <= '0';
partial_product_13(398) <= '0';
partial_product_13(399) <= '0';
partial_product_13(400) <= '0';
partial_product_13(401) <= '0';
partial_product_13(402) <= '0';
partial_product_13(403) <= '0';
partial_product_13(404) <= '0';
partial_product_13(405) <= '0';
partial_product_13(406) <= '0';
partial_product_13(407) <= '0';
partial_product_13(408) <= '0';
partial_product_13(409) <= '0';
partial_product_13(410) <= '0';
partial_product_13(411) <= '0';
partial_product_13(412) <= '0';
partial_product_13(413) <= '0';
partial_product_13(414) <= '0';
partial_product_13(415) <= '0';
partial_product_13(416) <= '0';
partial_product_13(417) <= '0';
partial_product_13(418) <= '0';
partial_product_13(419) <= '0';
partial_product_13(420) <= '0';
partial_product_13(421) <= '0';
partial_product_13(422) <= '0';
partial_product_13(423) <= '0';
partial_product_13(424) <= '0';
partial_product_13(425) <= '0';
partial_product_13(426) <= '0';
partial_product_13(427) <= '0';
partial_product_13(428) <= '0';
partial_product_13(429) <= '0';
partial_product_13(430) <= '0';
partial_product_13(431) <= '0';
partial_product_13(432) <= '0';
partial_product_13(433) <= '0';
partial_product_13(434) <= '0';
partial_product_13(435) <= '0';
partial_product_13(436) <= '0';
partial_product_13(437) <= '0';
partial_product_13(438) <= '0';
partial_product_13(439) <= '0';
partial_product_13(440) <= '0';
partial_product_13(441) <= '0';
partial_product_13(442) <= '0';
partial_product_13(443) <= '0';
partial_product_13(444) <= '0';
partial_product_13(445) <= '0';
partial_product_13(446) <= '0';
partial_product_13(447) <= '0';
partial_product_13(448) <= '0';
partial_product_13(449) <= '0';
partial_product_13(450) <= '0';
partial_product_13(451) <= '0';
partial_product_13(452) <= '0';
partial_product_13(453) <= '0';
partial_product_13(454) <= '0';
partial_product_13(455) <= '0';
partial_product_13(456) <= '0';
partial_product_13(457) <= '0';
partial_product_13(458) <= '0';
partial_product_13(459) <= '0';
partial_product_13(460) <= '0';
partial_product_13(461) <= '0';
partial_product_13(462) <= '0';
partial_product_13(463) <= '0';
partial_product_13(464) <= '0';
partial_product_13(465) <= '0';
partial_product_13(466) <= '0';
partial_product_13(467) <= '0';
partial_product_13(468) <= '0';
partial_product_13(469) <= '0';
partial_product_13(470) <= '0';
partial_product_13(471) <= '0';
partial_product_13(472) <= '0';
partial_product_13(473) <= '0';
partial_product_13(474) <= '0';
partial_product_13(475) <= '0';
partial_product_13(476) <= '0';
partial_product_13(477) <= '0';
partial_product_13(478) <= '0';
partial_product_13(479) <= '0';
partial_product_13(480) <= '0';
partial_product_13(481) <= '0';
partial_product_13(482) <= '0';
partial_product_13(483) <= '0';
partial_product_13(484) <= '0';
partial_product_13(485) <= '0';
partial_product_13(486) <= '0';
partial_product_13(487) <= '0';
partial_product_13(488) <= '0';
partial_product_13(489) <= '0';
partial_product_13(490) <= '0';
partial_product_13(491) <= '0';
partial_product_13(492) <= '0';
partial_product_13(493) <= '0';
partial_product_13(494) <= '0';
partial_product_13(495) <= '0';
partial_product_13(496) <= '0';
partial_product_13(497) <= '0';
partial_product_13(498) <= '0';
partial_product_13(499) <= '0';
partial_product_13(500) <= '0';
partial_product_13(501) <= '0';
partial_product_13(502) <= '0';
partial_product_13(503) <= '0';
partial_product_13(504) <= '0';
partial_product_13(505) <= '0';
partial_product_13(506) <= '0';
partial_product_13(507) <= '0';
partial_product_13(508) <= '0';
partial_product_13(509) <= '0';
partial_product_13(510) <= '0';
partial_product_13(511) <= '0';
partial_product_13(512) <= '0';
partial_product_14(0) <= '0';
partial_product_14(1) <= '0';
partial_product_14(2) <= '0';
partial_product_14(3) <= '0';
partial_product_14(4) <= '0';
partial_product_14(5) <= '0';
partial_product_14(6) <= '0';
partial_product_14(7) <= '0';
partial_product_14(8) <= '0';
partial_product_14(9) <= '0';
partial_product_14(10) <= '0';
partial_product_14(11) <= '0';
partial_product_14(12) <= '0';
partial_product_14(13) <= '0';
partial_product_14(14) <= '0';
partial_product_14(15) <= '0';
partial_product_14(16) <= '0';
partial_product_14(17) <= '0';
partial_product_14(18) <= '0';
partial_product_14(19) <= '0';
partial_product_14(20) <= '0';
partial_product_14(21) <= '0';
partial_product_14(22) <= '0';
partial_product_14(23) <= '0';
partial_product_14(24) <= '0';
partial_product_14(25) <= '0';
partial_product_14(26) <= '0';
partial_product_14(27) <= '0';
partial_product_14(28) <= '0';
partial_product_14(29) <= '0';
partial_product_14(30) <= '0';
partial_product_14(31) <= '0';
partial_product_14(32) <= '0';
partial_product_14(33) <= '0';
partial_product_14(34) <= '0';
partial_product_14(35) <= '0';
partial_product_14(36) <= '0';
partial_product_14(37) <= '0';
partial_product_14(38) <= '0';
partial_product_14(39) <= '0';
partial_product_14(40) <= '0';
partial_product_14(41) <= '0';
partial_product_14(42) <= '0';
partial_product_14(43) <= '0';
partial_product_14(44) <= '0';
partial_product_14(45) <= '0';
partial_product_14(46) <= '0';
partial_product_14(47) <= '0';
partial_product_14(48) <= '0';
partial_product_14(49) <= '0';
partial_product_14(50) <= '0';
partial_product_14(51) <= '0';
partial_product_14(52) <= '0';
partial_product_14(53) <= '0';
partial_product_14(54) <= '0';
partial_product_14(55) <= '0';
partial_product_14(56) <= '0';
partial_product_14(57) <= '0';
partial_product_14(58) <= '0';
partial_product_14(59) <= '0';
partial_product_14(60) <= '0';
partial_product_14(61) <= '0';
partial_product_14(62) <= '0';
partial_product_14(63) <= '0';
partial_product_14(64) <= '0';
partial_product_14(65) <= '0';
partial_product_14(66) <= '0';
partial_product_14(67) <= '0';
partial_product_14(68) <= '0';
partial_product_14(69) <= '0';
partial_product_14(70) <= '0';
partial_product_14(71) <= '0';
partial_product_14(72) <= '0';
partial_product_14(73) <= '0';
partial_product_14(74) <= '0';
partial_product_14(75) <= '0';
partial_product_14(76) <= '0';
partial_product_14(77) <= '0';
partial_product_14(78) <= '0';
partial_product_14(79) <= '0';
partial_product_14(80) <= '0';
partial_product_14(81) <= '0';
partial_product_14(82) <= '0';
partial_product_14(83) <= '0';
partial_product_14(84) <= '0';
partial_product_14(85) <= '0';
partial_product_14(86) <= '0';
partial_product_14(87) <= '0';
partial_product_14(88) <= '0';
partial_product_14(89) <= '0';
partial_product_14(90) <= '0';
partial_product_14(91) <= '0';
partial_product_14(92) <= '0';
partial_product_14(93) <= '0';
partial_product_14(94) <= '0';
partial_product_14(95) <= '0';
partial_product_14(96) <= '0';
partial_product_14(97) <= '0';
partial_product_14(98) <= '0';
partial_product_14(99) <= '0';
partial_product_14(100) <= '0';
partial_product_14(101) <= '0';
partial_product_14(102) <= '0';
partial_product_14(103) <= '0';
partial_product_14(104) <= '0';
partial_product_14(105) <= '0';
partial_product_14(106) <= '0';
partial_product_14(107) <= '0';
partial_product_14(108) <= '0';
partial_product_14(109) <= '0';
partial_product_14(110) <= '0';
partial_product_14(111) <= '0';
partial_product_14(112) <= '0';
partial_product_14(113) <= '0';
partial_product_14(114) <= '0';
partial_product_14(115) <= '0';
partial_product_14(116) <= '0';
partial_product_14(117) <= '0';
partial_product_14(118) <= '0';
partial_product_14(119) <= '0';
partial_product_14(120) <= '0';
partial_product_14(121) <= '0';
partial_product_14(122) <= '0';
partial_product_14(123) <= '0';
partial_product_14(124) <= '0';
partial_product_14(125) <= '0';
partial_product_14(126) <= '0';
partial_product_14(127) <= '0';
partial_product_14(128) <= '0';
partial_product_14(129) <= '0';
partial_product_14(130) <= '0';
partial_product_14(131) <= '0';
partial_product_14(132) <= '0';
partial_product_14(133) <= '0';
partial_product_14(134) <= '0';
partial_product_14(135) <= '0';
partial_product_14(136) <= '0';
partial_product_14(137) <= '0';
partial_product_14(138) <= '0';
partial_product_14(139) <= '0';
partial_product_14(140) <= '0';
partial_product_14(141) <= '0';
partial_product_14(142) <= '0';
partial_product_14(143) <= '0';
partial_product_14(144) <= temp_mult_48(144);
partial_product_14(145) <= temp_mult_48(145);
partial_product_14(146) <= temp_mult_48(146);
partial_product_14(147) <= temp_mult_48(147);
partial_product_14(148) <= temp_mult_48(148);
partial_product_14(149) <= temp_mult_48(149);
partial_product_14(150) <= temp_mult_48(150);
partial_product_14(151) <= temp_mult_48(151);
partial_product_14(152) <= temp_mult_48(152);
partial_product_14(153) <= temp_mult_48(153);
partial_product_14(154) <= temp_mult_48(154);
partial_product_14(155) <= temp_mult_48(155);
partial_product_14(156) <= temp_mult_48(156);
partial_product_14(157) <= temp_mult_48(157);
partial_product_14(158) <= temp_mult_48(158);
partial_product_14(159) <= temp_mult_48(159);
partial_product_14(160) <= temp_mult_48(160);
partial_product_14(161) <= temp_mult_48(161);
partial_product_14(162) <= temp_mult_48(162);
partial_product_14(163) <= temp_mult_48(163);
partial_product_14(164) <= temp_mult_48(164);
partial_product_14(165) <= temp_mult_48(165);
partial_product_14(166) <= temp_mult_48(166);
partial_product_14(167) <= temp_mult_48(167);
partial_product_14(168) <= temp_mult_48(168);
partial_product_14(169) <= temp_mult_48(169);
partial_product_14(170) <= temp_mult_48(170);
partial_product_14(171) <= temp_mult_48(171);
partial_product_14(172) <= temp_mult_48(172);
partial_product_14(173) <= temp_mult_48(173);
partial_product_14(174) <= temp_mult_48(174);
partial_product_14(175) <= temp_mult_48(175);
partial_product_14(176) <= temp_mult_48(176);
partial_product_14(177) <= temp_mult_48(177);
partial_product_14(178) <= temp_mult_48(178);
partial_product_14(179) <= temp_mult_48(179);
partial_product_14(180) <= temp_mult_48(180);
partial_product_14(181) <= temp_mult_48(181);
partial_product_14(182) <= temp_mult_48(182);
partial_product_14(183) <= temp_mult_48(183);
partial_product_14(184) <= temp_mult_48(184);
partial_product_14(185) <= temp_mult_57(185);
partial_product_14(186) <= temp_mult_57(186);
partial_product_14(187) <= temp_mult_57(187);
partial_product_14(188) <= temp_mult_57(188);
partial_product_14(189) <= temp_mult_57(189);
partial_product_14(190) <= temp_mult_57(190);
partial_product_14(191) <= temp_mult_57(191);
partial_product_14(192) <= temp_mult_57(192);
partial_product_14(193) <= temp_mult_57(193);
partial_product_14(194) <= temp_mult_57(194);
partial_product_14(195) <= temp_mult_57(195);
partial_product_14(196) <= temp_mult_57(196);
partial_product_14(197) <= temp_mult_57(197);
partial_product_14(198) <= temp_mult_57(198);
partial_product_14(199) <= temp_mult_57(199);
partial_product_14(200) <= temp_mult_57(200);
partial_product_14(201) <= temp_mult_57(201);
partial_product_14(202) <= temp_mult_57(202);
partial_product_14(203) <= temp_mult_57(203);
partial_product_14(204) <= temp_mult_57(204);
partial_product_14(205) <= temp_mult_57(205);
partial_product_14(206) <= temp_mult_57(206);
partial_product_14(207) <= temp_mult_57(207);
partial_product_14(208) <= temp_mult_57(208);
partial_product_14(209) <= temp_mult_57(209);
partial_product_14(210) <= temp_mult_57(210);
partial_product_14(211) <= temp_mult_57(211);
partial_product_14(212) <= temp_mult_57(212);
partial_product_14(213) <= temp_mult_57(213);
partial_product_14(214) <= temp_mult_57(214);
partial_product_14(215) <= temp_mult_57(215);
partial_product_14(216) <= temp_mult_57(216);
partial_product_14(217) <= temp_mult_57(217);
partial_product_14(218) <= temp_mult_57(218);
partial_product_14(219) <= temp_mult_57(219);
partial_product_14(220) <= temp_mult_57(220);
partial_product_14(221) <= temp_mult_57(221);
partial_product_14(222) <= temp_mult_57(222);
partial_product_14(223) <= temp_mult_57(223);
partial_product_14(224) <= temp_mult_57(224);
partial_product_14(225) <= temp_mult_57(225);
partial_product_14(226) <= temp_mult_66(226);
partial_product_14(227) <= temp_mult_66(227);
partial_product_14(228) <= temp_mult_66(228);
partial_product_14(229) <= temp_mult_66(229);
partial_product_14(230) <= temp_mult_66(230);
partial_product_14(231) <= temp_mult_66(231);
partial_product_14(232) <= temp_mult_66(232);
partial_product_14(233) <= temp_mult_66(233);
partial_product_14(234) <= temp_mult_66(234);
partial_product_14(235) <= temp_mult_66(235);
partial_product_14(236) <= temp_mult_66(236);
partial_product_14(237) <= temp_mult_66(237);
partial_product_14(238) <= temp_mult_66(238);
partial_product_14(239) <= temp_mult_66(239);
partial_product_14(240) <= temp_mult_66(240);
partial_product_14(241) <= temp_mult_66(241);
partial_product_14(242) <= temp_mult_66(242);
partial_product_14(243) <= temp_mult_66(243);
partial_product_14(244) <= temp_mult_66(244);
partial_product_14(245) <= temp_mult_66(245);
partial_product_14(246) <= temp_mult_66(246);
partial_product_14(247) <= temp_mult_66(247);
partial_product_14(248) <= temp_mult_66(248);
partial_product_14(249) <= temp_mult_66(249);
partial_product_14(250) <= temp_mult_66(250);
partial_product_14(251) <= temp_mult_66(251);
partial_product_14(252) <= temp_mult_66(252);
partial_product_14(253) <= temp_mult_66(253);
partial_product_14(254) <= temp_mult_66(254);
partial_product_14(255) <= temp_mult_66(255);
partial_product_14(256) <= temp_mult_66(256);
partial_product_14(257) <= temp_mult_66(257);
partial_product_14(258) <= temp_mult_66(258);
partial_product_14(259) <= temp_mult_66(259);
partial_product_14(260) <= temp_mult_66(260);
partial_product_14(261) <= temp_mult_66(261);
partial_product_14(262) <= temp_mult_66(262);
partial_product_14(263) <= temp_mult_66(263);
partial_product_14(264) <= temp_mult_66(264);
partial_product_14(265) <= temp_mult_66(265);
partial_product_14(266) <= temp_mult_66(266);
partial_product_14(267) <= temp_mult_75(267);
partial_product_14(268) <= temp_mult_75(268);
partial_product_14(269) <= temp_mult_75(269);
partial_product_14(270) <= temp_mult_75(270);
partial_product_14(271) <= temp_mult_75(271);
partial_product_14(272) <= temp_mult_75(272);
partial_product_14(273) <= temp_mult_75(273);
partial_product_14(274) <= temp_mult_75(274);
partial_product_14(275) <= temp_mult_75(275);
partial_product_14(276) <= temp_mult_75(276);
partial_product_14(277) <= temp_mult_75(277);
partial_product_14(278) <= temp_mult_75(278);
partial_product_14(279) <= temp_mult_75(279);
partial_product_14(280) <= temp_mult_75(280);
partial_product_14(281) <= temp_mult_75(281);
partial_product_14(282) <= temp_mult_75(282);
partial_product_14(283) <= temp_mult_75(283);
partial_product_14(284) <= temp_mult_75(284);
partial_product_14(285) <= temp_mult_75(285);
partial_product_14(286) <= temp_mult_75(286);
partial_product_14(287) <= temp_mult_75(287);
partial_product_14(288) <= temp_mult_75(288);
partial_product_14(289) <= temp_mult_75(289);
partial_product_14(290) <= temp_mult_75(290);
partial_product_14(291) <= temp_mult_75(291);
partial_product_14(292) <= temp_mult_75(292);
partial_product_14(293) <= temp_mult_75(293);
partial_product_14(294) <= temp_mult_75(294);
partial_product_14(295) <= temp_mult_75(295);
partial_product_14(296) <= temp_mult_75(296);
partial_product_14(297) <= temp_mult_75(297);
partial_product_14(298) <= temp_mult_75(298);
partial_product_14(299) <= temp_mult_75(299);
partial_product_14(300) <= temp_mult_75(300);
partial_product_14(301) <= temp_mult_75(301);
partial_product_14(302) <= temp_mult_75(302);
partial_product_14(303) <= temp_mult_75(303);
partial_product_14(304) <= temp_mult_75(304);
partial_product_14(305) <= temp_mult_75(305);
partial_product_14(306) <= temp_mult_75(306);
partial_product_14(307) <= temp_mult_75(307);
partial_product_14(308) <= '0';
partial_product_14(309) <= '0';
partial_product_14(310) <= temp_mult_110(310);
partial_product_14(311) <= temp_mult_110(311);
partial_product_14(312) <= temp_mult_110(312);
partial_product_14(313) <= temp_mult_110(313);
partial_product_14(314) <= temp_mult_110(314);
partial_product_14(315) <= temp_mult_110(315);
partial_product_14(316) <= temp_mult_110(316);
partial_product_14(317) <= temp_mult_110(317);
partial_product_14(318) <= temp_mult_110(318);
partial_product_14(319) <= temp_mult_110(319);
partial_product_14(320) <= temp_mult_110(320);
partial_product_14(321) <= temp_mult_110(321);
partial_product_14(322) <= temp_mult_110(322);
partial_product_14(323) <= temp_mult_110(323);
partial_product_14(324) <= temp_mult_110(324);
partial_product_14(325) <= temp_mult_110(325);
partial_product_14(326) <= temp_mult_110(326);
partial_product_14(327) <= temp_mult_110(327);
partial_product_14(328) <= temp_mult_110(328);
partial_product_14(329) <= temp_mult_110(329);
partial_product_14(330) <= temp_mult_110(330);
partial_product_14(331) <= temp_mult_110(331);
partial_product_14(332) <= temp_mult_110(332);
partial_product_14(333) <= temp_mult_110(333);
partial_product_14(334) <= temp_mult_110(334);
partial_product_14(335) <= temp_mult_110(335);
partial_product_14(336) <= temp_mult_110(336);
partial_product_14(337) <= temp_mult_110(337);
partial_product_14(338) <= temp_mult_110(338);
partial_product_14(339) <= temp_mult_110(339);
partial_product_14(340) <= temp_mult_110(340);
partial_product_14(341) <= temp_mult_110(341);
partial_product_14(342) <= temp_mult_110(342);
partial_product_14(343) <= temp_mult_110(343);
partial_product_14(344) <= temp_mult_110(344);
partial_product_14(345) <= temp_mult_110(345);
partial_product_14(346) <= temp_mult_110(346);
partial_product_14(347) <= temp_mult_110(347);
partial_product_14(348) <= temp_mult_110(348);
partial_product_14(349) <= temp_mult_110(349);
partial_product_14(350) <= temp_mult_110(350);
partial_product_14(351) <= '0';
partial_product_14(352) <= '0';
partial_product_14(353) <= '0';
partial_product_14(354) <= '0';
partial_product_14(355) <= '0';
partial_product_14(356) <= '0';
partial_product_14(357) <= '0';
partial_product_14(358) <= temp_mult_150(358);
partial_product_14(359) <= temp_mult_150(359);
partial_product_14(360) <= temp_mult_150(360);
partial_product_14(361) <= temp_mult_150(361);
partial_product_14(362) <= temp_mult_150(362);
partial_product_14(363) <= temp_mult_150(363);
partial_product_14(364) <= temp_mult_150(364);
partial_product_14(365) <= temp_mult_150(365);
partial_product_14(366) <= temp_mult_150(366);
partial_product_14(367) <= temp_mult_150(367);
partial_product_14(368) <= temp_mult_150(368);
partial_product_14(369) <= temp_mult_150(369);
partial_product_14(370) <= temp_mult_150(370);
partial_product_14(371) <= temp_mult_150(371);
partial_product_14(372) <= temp_mult_150(372);
partial_product_14(373) <= temp_mult_150(373);
partial_product_14(374) <= temp_mult_150(374);
partial_product_14(375) <= temp_mult_150(375);
partial_product_14(376) <= temp_mult_150(376);
partial_product_14(377) <= temp_mult_150(377);
partial_product_14(378) <= temp_mult_150(378);
partial_product_14(379) <= temp_mult_150(379);
partial_product_14(380) <= temp_mult_150(380);
partial_product_14(381) <= temp_mult_150(381);
partial_product_14(382) <= temp_mult_150(382);
partial_product_14(383) <= temp_mult_150(383);
partial_product_14(384) <= temp_mult_150(384);
partial_product_14(385) <= temp_mult_150(385);
partial_product_14(386) <= temp_mult_150(386);
partial_product_14(387) <= temp_mult_150(387);
partial_product_14(388) <= temp_mult_150(388);
partial_product_14(389) <= temp_mult_150(389);
partial_product_14(390) <= temp_mult_150(390);
partial_product_14(391) <= temp_mult_150(391);
partial_product_14(392) <= temp_mult_150(392);
partial_product_14(393) <= temp_mult_150(393);
partial_product_14(394) <= temp_mult_150(394);
partial_product_14(395) <= temp_mult_150(395);
partial_product_14(396) <= temp_mult_150(396);
partial_product_14(397) <= temp_mult_150(397);
partial_product_14(398) <= temp_mult_150(398);
partial_product_14(399) <= '0';
partial_product_14(400) <= '0';
partial_product_14(401) <= '0';
partial_product_14(402) <= '0';
partial_product_14(403) <= '0';
partial_product_14(404) <= '0';
partial_product_14(405) <= '0';
partial_product_14(406) <= '0';
partial_product_14(407) <= '0';
partial_product_14(408) <= '0';
partial_product_14(409) <= '0';
partial_product_14(410) <= '0';
partial_product_14(411) <= '0';
partial_product_14(412) <= '0';
partial_product_14(413) <= '0';
partial_product_14(414) <= '0';
partial_product_14(415) <= '0';
partial_product_14(416) <= '0';
partial_product_14(417) <= '0';
partial_product_14(418) <= '0';
partial_product_14(419) <= '0';
partial_product_14(420) <= '0';
partial_product_14(421) <= '0';
partial_product_14(422) <= '0';
partial_product_14(423) <= '0';
partial_product_14(424) <= '0';
partial_product_14(425) <= '0';
partial_product_14(426) <= '0';
partial_product_14(427) <= '0';
partial_product_14(428) <= '0';
partial_product_14(429) <= '0';
partial_product_14(430) <= '0';
partial_product_14(431) <= '0';
partial_product_14(432) <= '0';
partial_product_14(433) <= '0';
partial_product_14(434) <= '0';
partial_product_14(435) <= '0';
partial_product_14(436) <= '0';
partial_product_14(437) <= '0';
partial_product_14(438) <= '0';
partial_product_14(439) <= '0';
partial_product_14(440) <= '0';
partial_product_14(441) <= '0';
partial_product_14(442) <= '0';
partial_product_14(443) <= '0';
partial_product_14(444) <= '0';
partial_product_14(445) <= '0';
partial_product_14(446) <= '0';
partial_product_14(447) <= '0';
partial_product_14(448) <= '0';
partial_product_14(449) <= '0';
partial_product_14(450) <= '0';
partial_product_14(451) <= '0';
partial_product_14(452) <= '0';
partial_product_14(453) <= '0';
partial_product_14(454) <= '0';
partial_product_14(455) <= '0';
partial_product_14(456) <= '0';
partial_product_14(457) <= '0';
partial_product_14(458) <= '0';
partial_product_14(459) <= '0';
partial_product_14(460) <= '0';
partial_product_14(461) <= '0';
partial_product_14(462) <= '0';
partial_product_14(463) <= '0';
partial_product_14(464) <= '0';
partial_product_14(465) <= '0';
partial_product_14(466) <= '0';
partial_product_14(467) <= '0';
partial_product_14(468) <= '0';
partial_product_14(469) <= '0';
partial_product_14(470) <= '0';
partial_product_14(471) <= '0';
partial_product_14(472) <= '0';
partial_product_14(473) <= '0';
partial_product_14(474) <= '0';
partial_product_14(475) <= '0';
partial_product_14(476) <= '0';
partial_product_14(477) <= '0';
partial_product_14(478) <= '0';
partial_product_14(479) <= '0';
partial_product_14(480) <= '0';
partial_product_14(481) <= '0';
partial_product_14(482) <= '0';
partial_product_14(483) <= '0';
partial_product_14(484) <= '0';
partial_product_14(485) <= '0';
partial_product_14(486) <= '0';
partial_product_14(487) <= '0';
partial_product_14(488) <= '0';
partial_product_14(489) <= '0';
partial_product_14(490) <= '0';
partial_product_14(491) <= '0';
partial_product_14(492) <= '0';
partial_product_14(493) <= '0';
partial_product_14(494) <= '0';
partial_product_14(495) <= '0';
partial_product_14(496) <= '0';
partial_product_14(497) <= '0';
partial_product_14(498) <= '0';
partial_product_14(499) <= '0';
partial_product_14(500) <= '0';
partial_product_14(501) <= '0';
partial_product_14(502) <= '0';
partial_product_14(503) <= '0';
partial_product_14(504) <= '0';
partial_product_14(505) <= '0';
partial_product_14(506) <= '0';
partial_product_14(507) <= '0';
partial_product_14(508) <= '0';
partial_product_14(509) <= '0';
partial_product_14(510) <= '0';
partial_product_14(511) <= '0';
partial_product_14(512) <= '0';
partial_product_15(0) <= '0';
partial_product_15(1) <= '0';
partial_product_15(2) <= '0';
partial_product_15(3) <= '0';
partial_product_15(4) <= '0';
partial_product_15(5) <= '0';
partial_product_15(6) <= '0';
partial_product_15(7) <= '0';
partial_product_15(8) <= '0';
partial_product_15(9) <= '0';
partial_product_15(10) <= '0';
partial_product_15(11) <= '0';
partial_product_15(12) <= '0';
partial_product_15(13) <= '0';
partial_product_15(14) <= '0';
partial_product_15(15) <= '0';
partial_product_15(16) <= '0';
partial_product_15(17) <= '0';
partial_product_15(18) <= '0';
partial_product_15(19) <= '0';
partial_product_15(20) <= '0';
partial_product_15(21) <= '0';
partial_product_15(22) <= '0';
partial_product_15(23) <= '0';
partial_product_15(24) <= '0';
partial_product_15(25) <= '0';
partial_product_15(26) <= '0';
partial_product_15(27) <= '0';
partial_product_15(28) <= '0';
partial_product_15(29) <= '0';
partial_product_15(30) <= '0';
partial_product_15(31) <= '0';
partial_product_15(32) <= '0';
partial_product_15(33) <= '0';
partial_product_15(34) <= '0';
partial_product_15(35) <= '0';
partial_product_15(36) <= '0';
partial_product_15(37) <= '0';
partial_product_15(38) <= '0';
partial_product_15(39) <= '0';
partial_product_15(40) <= '0';
partial_product_15(41) <= '0';
partial_product_15(42) <= '0';
partial_product_15(43) <= '0';
partial_product_15(44) <= '0';
partial_product_15(45) <= '0';
partial_product_15(46) <= '0';
partial_product_15(47) <= '0';
partial_product_15(48) <= '0';
partial_product_15(49) <= '0';
partial_product_15(50) <= '0';
partial_product_15(51) <= '0';
partial_product_15(52) <= '0';
partial_product_15(53) <= '0';
partial_product_15(54) <= '0';
partial_product_15(55) <= '0';
partial_product_15(56) <= '0';
partial_product_15(57) <= '0';
partial_product_15(58) <= '0';
partial_product_15(59) <= '0';
partial_product_15(60) <= '0';
partial_product_15(61) <= '0';
partial_product_15(62) <= '0';
partial_product_15(63) <= '0';
partial_product_15(64) <= '0';
partial_product_15(65) <= '0';
partial_product_15(66) <= '0';
partial_product_15(67) <= '0';
partial_product_15(68) <= '0';
partial_product_15(69) <= '0';
partial_product_15(70) <= '0';
partial_product_15(71) <= '0';
partial_product_15(72) <= '0';
partial_product_15(73) <= '0';
partial_product_15(74) <= '0';
partial_product_15(75) <= '0';
partial_product_15(76) <= '0';
partial_product_15(77) <= '0';
partial_product_15(78) <= '0';
partial_product_15(79) <= '0';
partial_product_15(80) <= '0';
partial_product_15(81) <= '0';
partial_product_15(82) <= '0';
partial_product_15(83) <= '0';
partial_product_15(84) <= '0';
partial_product_15(85) <= '0';
partial_product_15(86) <= '0';
partial_product_15(87) <= '0';
partial_product_15(88) <= '0';
partial_product_15(89) <= '0';
partial_product_15(90) <= '0';
partial_product_15(91) <= '0';
partial_product_15(92) <= '0';
partial_product_15(93) <= '0';
partial_product_15(94) <= '0';
partial_product_15(95) <= '0';
partial_product_15(96) <= '0';
partial_product_15(97) <= '0';
partial_product_15(98) <= '0';
partial_product_15(99) <= '0';
partial_product_15(100) <= '0';
partial_product_15(101) <= '0';
partial_product_15(102) <= '0';
partial_product_15(103) <= '0';
partial_product_15(104) <= '0';
partial_product_15(105) <= '0';
partial_product_15(106) <= '0';
partial_product_15(107) <= '0';
partial_product_15(108) <= '0';
partial_product_15(109) <= '0';
partial_product_15(110) <= '0';
partial_product_15(111) <= '0';
partial_product_15(112) <= '0';
partial_product_15(113) <= '0';
partial_product_15(114) <= '0';
partial_product_15(115) <= '0';
partial_product_15(116) <= '0';
partial_product_15(117) <= '0';
partial_product_15(118) <= '0';
partial_product_15(119) <= '0';
partial_product_15(120) <= '0';
partial_product_15(121) <= '0';
partial_product_15(122) <= '0';
partial_product_15(123) <= '0';
partial_product_15(124) <= '0';
partial_product_15(125) <= '0';
partial_product_15(126) <= '0';
partial_product_15(127) <= '0';
partial_product_15(128) <= '0';
partial_product_15(129) <= '0';
partial_product_15(130) <= '0';
partial_product_15(131) <= '0';
partial_product_15(132) <= '0';
partial_product_15(133) <= '0';
partial_product_15(134) <= '0';
partial_product_15(135) <= '0';
partial_product_15(136) <= '0';
partial_product_15(137) <= '0';
partial_product_15(138) <= '0';
partial_product_15(139) <= '0';
partial_product_15(140) <= '0';
partial_product_15(141) <= '0';
partial_product_15(142) <= '0';
partial_product_15(143) <= '0';
partial_product_15(144) <= '0';
partial_product_15(145) <= '0';
partial_product_15(146) <= '0';
partial_product_15(147) <= '0';
partial_product_15(148) <= '0';
partial_product_15(149) <= '0';
partial_product_15(150) <= '0';
partial_product_15(151) <= '0';
partial_product_15(152) <= '0';
partial_product_15(153) <= temp_mult_81(153);
partial_product_15(154) <= temp_mult_81(154);
partial_product_15(155) <= temp_mult_81(155);
partial_product_15(156) <= temp_mult_81(156);
partial_product_15(157) <= temp_mult_81(157);
partial_product_15(158) <= temp_mult_81(158);
partial_product_15(159) <= temp_mult_81(159);
partial_product_15(160) <= temp_mult_81(160);
partial_product_15(161) <= temp_mult_81(161);
partial_product_15(162) <= temp_mult_81(162);
partial_product_15(163) <= temp_mult_81(163);
partial_product_15(164) <= temp_mult_81(164);
partial_product_15(165) <= temp_mult_81(165);
partial_product_15(166) <= temp_mult_81(166);
partial_product_15(167) <= temp_mult_81(167);
partial_product_15(168) <= temp_mult_81(168);
partial_product_15(169) <= temp_mult_81(169);
partial_product_15(170) <= temp_mult_81(170);
partial_product_15(171) <= temp_mult_81(171);
partial_product_15(172) <= temp_mult_81(172);
partial_product_15(173) <= temp_mult_81(173);
partial_product_15(174) <= temp_mult_81(174);
partial_product_15(175) <= temp_mult_81(175);
partial_product_15(176) <= temp_mult_81(176);
partial_product_15(177) <= temp_mult_81(177);
partial_product_15(178) <= temp_mult_81(178);
partial_product_15(179) <= temp_mult_81(179);
partial_product_15(180) <= temp_mult_81(180);
partial_product_15(181) <= temp_mult_81(181);
partial_product_15(182) <= temp_mult_81(182);
partial_product_15(183) <= temp_mult_81(183);
partial_product_15(184) <= temp_mult_81(184);
partial_product_15(185) <= temp_mult_81(185);
partial_product_15(186) <= temp_mult_81(186);
partial_product_15(187) <= temp_mult_81(187);
partial_product_15(188) <= temp_mult_81(188);
partial_product_15(189) <= temp_mult_81(189);
partial_product_15(190) <= temp_mult_81(190);
partial_product_15(191) <= temp_mult_81(191);
partial_product_15(192) <= temp_mult_81(192);
partial_product_15(193) <= temp_mult_81(193);
partial_product_15(194) <= temp_mult_90(194);
partial_product_15(195) <= temp_mult_90(195);
partial_product_15(196) <= temp_mult_90(196);
partial_product_15(197) <= temp_mult_90(197);
partial_product_15(198) <= temp_mult_90(198);
partial_product_15(199) <= temp_mult_90(199);
partial_product_15(200) <= temp_mult_90(200);
partial_product_15(201) <= temp_mult_90(201);
partial_product_15(202) <= temp_mult_90(202);
partial_product_15(203) <= temp_mult_90(203);
partial_product_15(204) <= temp_mult_90(204);
partial_product_15(205) <= temp_mult_90(205);
partial_product_15(206) <= temp_mult_90(206);
partial_product_15(207) <= temp_mult_90(207);
partial_product_15(208) <= temp_mult_90(208);
partial_product_15(209) <= temp_mult_90(209);
partial_product_15(210) <= temp_mult_90(210);
partial_product_15(211) <= temp_mult_90(211);
partial_product_15(212) <= temp_mult_90(212);
partial_product_15(213) <= temp_mult_90(213);
partial_product_15(214) <= temp_mult_90(214);
partial_product_15(215) <= temp_mult_90(215);
partial_product_15(216) <= temp_mult_90(216);
partial_product_15(217) <= temp_mult_90(217);
partial_product_15(218) <= temp_mult_90(218);
partial_product_15(219) <= temp_mult_90(219);
partial_product_15(220) <= temp_mult_90(220);
partial_product_15(221) <= temp_mult_90(221);
partial_product_15(222) <= temp_mult_90(222);
partial_product_15(223) <= temp_mult_90(223);
partial_product_15(224) <= temp_mult_90(224);
partial_product_15(225) <= temp_mult_90(225);
partial_product_15(226) <= temp_mult_90(226);
partial_product_15(227) <= temp_mult_90(227);
partial_product_15(228) <= temp_mult_90(228);
partial_product_15(229) <= temp_mult_90(229);
partial_product_15(230) <= temp_mult_90(230);
partial_product_15(231) <= temp_mult_90(231);
partial_product_15(232) <= temp_mult_90(232);
partial_product_15(233) <= temp_mult_90(233);
partial_product_15(234) <= temp_mult_90(234);
partial_product_15(235) <= temp_mult_99(235);
partial_product_15(236) <= temp_mult_99(236);
partial_product_15(237) <= temp_mult_99(237);
partial_product_15(238) <= temp_mult_99(238);
partial_product_15(239) <= temp_mult_99(239);
partial_product_15(240) <= temp_mult_99(240);
partial_product_15(241) <= temp_mult_99(241);
partial_product_15(242) <= temp_mult_99(242);
partial_product_15(243) <= temp_mult_99(243);
partial_product_15(244) <= temp_mult_99(244);
partial_product_15(245) <= temp_mult_99(245);
partial_product_15(246) <= temp_mult_99(246);
partial_product_15(247) <= temp_mult_99(247);
partial_product_15(248) <= temp_mult_99(248);
partial_product_15(249) <= temp_mult_99(249);
partial_product_15(250) <= temp_mult_99(250);
partial_product_15(251) <= temp_mult_99(251);
partial_product_15(252) <= temp_mult_99(252);
partial_product_15(253) <= temp_mult_99(253);
partial_product_15(254) <= temp_mult_99(254);
partial_product_15(255) <= temp_mult_99(255);
partial_product_15(256) <= temp_mult_99(256);
partial_product_15(257) <= temp_mult_99(257);
partial_product_15(258) <= temp_mult_99(258);
partial_product_15(259) <= temp_mult_99(259);
partial_product_15(260) <= temp_mult_99(260);
partial_product_15(261) <= temp_mult_99(261);
partial_product_15(262) <= temp_mult_99(262);
partial_product_15(263) <= temp_mult_99(263);
partial_product_15(264) <= temp_mult_99(264);
partial_product_15(265) <= temp_mult_99(265);
partial_product_15(266) <= temp_mult_99(266);
partial_product_15(267) <= temp_mult_99(267);
partial_product_15(268) <= temp_mult_99(268);
partial_product_15(269) <= temp_mult_99(269);
partial_product_15(270) <= temp_mult_99(270);
partial_product_15(271) <= temp_mult_99(271);
partial_product_15(272) <= temp_mult_99(272);
partial_product_15(273) <= temp_mult_99(273);
partial_product_15(274) <= temp_mult_99(274);
partial_product_15(275) <= temp_mult_99(275);
partial_product_15(276) <= temp_mult_108(276);
partial_product_15(277) <= temp_mult_108(277);
partial_product_15(278) <= temp_mult_108(278);
partial_product_15(279) <= temp_mult_108(279);
partial_product_15(280) <= temp_mult_108(280);
partial_product_15(281) <= temp_mult_108(281);
partial_product_15(282) <= temp_mult_108(282);
partial_product_15(283) <= temp_mult_108(283);
partial_product_15(284) <= temp_mult_108(284);
partial_product_15(285) <= temp_mult_108(285);
partial_product_15(286) <= temp_mult_108(286);
partial_product_15(287) <= temp_mult_108(287);
partial_product_15(288) <= temp_mult_108(288);
partial_product_15(289) <= temp_mult_108(289);
partial_product_15(290) <= temp_mult_108(290);
partial_product_15(291) <= temp_mult_108(291);
partial_product_15(292) <= temp_mult_108(292);
partial_product_15(293) <= temp_mult_108(293);
partial_product_15(294) <= temp_mult_108(294);
partial_product_15(295) <= temp_mult_108(295);
partial_product_15(296) <= temp_mult_108(296);
partial_product_15(297) <= temp_mult_108(297);
partial_product_15(298) <= temp_mult_108(298);
partial_product_15(299) <= temp_mult_108(299);
partial_product_15(300) <= temp_mult_108(300);
partial_product_15(301) <= temp_mult_108(301);
partial_product_15(302) <= temp_mult_108(302);
partial_product_15(303) <= temp_mult_108(303);
partial_product_15(304) <= temp_mult_108(304);
partial_product_15(305) <= temp_mult_108(305);
partial_product_15(306) <= temp_mult_108(306);
partial_product_15(307) <= temp_mult_108(307);
partial_product_15(308) <= temp_mult_108(308);
partial_product_15(309) <= temp_mult_108(309);
partial_product_15(310) <= temp_mult_108(310);
partial_product_15(311) <= temp_mult_108(311);
partial_product_15(312) <= temp_mult_108(312);
partial_product_15(313) <= temp_mult_108(313);
partial_product_15(314) <= temp_mult_108(314);
partial_product_15(315) <= temp_mult_108(315);
partial_product_15(316) <= temp_mult_108(316);
partial_product_15(317) <= temp_mult_117(317);
partial_product_15(318) <= temp_mult_117(318);
partial_product_15(319) <= temp_mult_117(319);
partial_product_15(320) <= temp_mult_117(320);
partial_product_15(321) <= temp_mult_117(321);
partial_product_15(322) <= temp_mult_117(322);
partial_product_15(323) <= temp_mult_117(323);
partial_product_15(324) <= temp_mult_117(324);
partial_product_15(325) <= temp_mult_117(325);
partial_product_15(326) <= temp_mult_117(326);
partial_product_15(327) <= temp_mult_117(327);
partial_product_15(328) <= temp_mult_117(328);
partial_product_15(329) <= temp_mult_117(329);
partial_product_15(330) <= temp_mult_117(330);
partial_product_15(331) <= temp_mult_117(331);
partial_product_15(332) <= temp_mult_117(332);
partial_product_15(333) <= temp_mult_117(333);
partial_product_15(334) <= temp_mult_117(334);
partial_product_15(335) <= temp_mult_117(335);
partial_product_15(336) <= temp_mult_117(336);
partial_product_15(337) <= temp_mult_117(337);
partial_product_15(338) <= temp_mult_117(338);
partial_product_15(339) <= temp_mult_117(339);
partial_product_15(340) <= temp_mult_117(340);
partial_product_15(341) <= temp_mult_117(341);
partial_product_15(342) <= temp_mult_117(342);
partial_product_15(343) <= temp_mult_117(343);
partial_product_15(344) <= temp_mult_117(344);
partial_product_15(345) <= temp_mult_117(345);
partial_product_15(346) <= temp_mult_117(346);
partial_product_15(347) <= temp_mult_117(347);
partial_product_15(348) <= temp_mult_117(348);
partial_product_15(349) <= temp_mult_117(349);
partial_product_15(350) <= temp_mult_117(350);
partial_product_15(351) <= temp_mult_117(351);
partial_product_15(352) <= temp_mult_117(352);
partial_product_15(353) <= temp_mult_117(353);
partial_product_15(354) <= temp_mult_117(354);
partial_product_15(355) <= temp_mult_117(355);
partial_product_15(356) <= temp_mult_117(356);
partial_product_15(357) <= temp_mult_117(357);
partial_product_15(358) <= '0';
partial_product_15(359) <= '0';
partial_product_15(360) <= '0';
partial_product_15(361) <= '0';
partial_product_15(362) <= '0';
partial_product_15(363) <= '0';
partial_product_15(364) <= '0';
partial_product_15(365) <= '0';
partial_product_15(366) <= '0';
partial_product_15(367) <= '0';
partial_product_15(368) <= '0';
partial_product_15(369) <= '0';
partial_product_15(370) <= '0';
partial_product_15(371) <= '0';
partial_product_15(372) <= '0';
partial_product_15(373) <= '0';
partial_product_15(374) <= '0';
partial_product_15(375) <= '0';
partial_product_15(376) <= '0';
partial_product_15(377) <= '0';
partial_product_15(378) <= '0';
partial_product_15(379) <= '0';
partial_product_15(380) <= '0';
partial_product_15(381) <= '0';
partial_product_15(382) <= '0';
partial_product_15(383) <= '0';
partial_product_15(384) <= '0';
partial_product_15(385) <= '0';
partial_product_15(386) <= '0';
partial_product_15(387) <= '0';
partial_product_15(388) <= '0';
partial_product_15(389) <= '0';
partial_product_15(390) <= '0';
partial_product_15(391) <= '0';
partial_product_15(392) <= '0';
partial_product_15(393) <= '0';
partial_product_15(394) <= '0';
partial_product_15(395) <= '0';
partial_product_15(396) <= '0';
partial_product_15(397) <= '0';
partial_product_15(398) <= '0';
partial_product_15(399) <= '0';
partial_product_15(400) <= '0';
partial_product_15(401) <= '0';
partial_product_15(402) <= '0';
partial_product_15(403) <= '0';
partial_product_15(404) <= '0';
partial_product_15(405) <= '0';
partial_product_15(406) <= '0';
partial_product_15(407) <= '0';
partial_product_15(408) <= '0';
partial_product_15(409) <= '0';
partial_product_15(410) <= '0';
partial_product_15(411) <= '0';
partial_product_15(412) <= '0';
partial_product_15(413) <= '0';
partial_product_15(414) <= '0';
partial_product_15(415) <= '0';
partial_product_15(416) <= '0';
partial_product_15(417) <= '0';
partial_product_15(418) <= '0';
partial_product_15(419) <= '0';
partial_product_15(420) <= '0';
partial_product_15(421) <= '0';
partial_product_15(422) <= '0';
partial_product_15(423) <= '0';
partial_product_15(424) <= '0';
partial_product_15(425) <= '0';
partial_product_15(426) <= '0';
partial_product_15(427) <= '0';
partial_product_15(428) <= '0';
partial_product_15(429) <= '0';
partial_product_15(430) <= '0';
partial_product_15(431) <= '0';
partial_product_15(432) <= '0';
partial_product_15(433) <= '0';
partial_product_15(434) <= '0';
partial_product_15(435) <= '0';
partial_product_15(436) <= '0';
partial_product_15(437) <= '0';
partial_product_15(438) <= '0';
partial_product_15(439) <= '0';
partial_product_15(440) <= '0';
partial_product_15(441) <= '0';
partial_product_15(442) <= '0';
partial_product_15(443) <= '0';
partial_product_15(444) <= '0';
partial_product_15(445) <= '0';
partial_product_15(446) <= '0';
partial_product_15(447) <= '0';
partial_product_15(448) <= '0';
partial_product_15(449) <= '0';
partial_product_15(450) <= '0';
partial_product_15(451) <= '0';
partial_product_15(452) <= '0';
partial_product_15(453) <= '0';
partial_product_15(454) <= '0';
partial_product_15(455) <= '0';
partial_product_15(456) <= '0';
partial_product_15(457) <= '0';
partial_product_15(458) <= '0';
partial_product_15(459) <= '0';
partial_product_15(460) <= '0';
partial_product_15(461) <= '0';
partial_product_15(462) <= '0';
partial_product_15(463) <= '0';
partial_product_15(464) <= '0';
partial_product_15(465) <= '0';
partial_product_15(466) <= '0';
partial_product_15(467) <= '0';
partial_product_15(468) <= '0';
partial_product_15(469) <= '0';
partial_product_15(470) <= '0';
partial_product_15(471) <= '0';
partial_product_15(472) <= '0';
partial_product_15(473) <= '0';
partial_product_15(474) <= '0';
partial_product_15(475) <= '0';
partial_product_15(476) <= '0';
partial_product_15(477) <= '0';
partial_product_15(478) <= '0';
partial_product_15(479) <= '0';
partial_product_15(480) <= '0';
partial_product_15(481) <= '0';
partial_product_15(482) <= '0';
partial_product_15(483) <= '0';
partial_product_15(484) <= '0';
partial_product_15(485) <= '0';
partial_product_15(486) <= '0';
partial_product_15(487) <= '0';
partial_product_15(488) <= '0';
partial_product_15(489) <= '0';
partial_product_15(490) <= '0';
partial_product_15(491) <= '0';
partial_product_15(492) <= '0';
partial_product_15(493) <= '0';
partial_product_15(494) <= '0';
partial_product_15(495) <= '0';
partial_product_15(496) <= '0';
partial_product_15(497) <= '0';
partial_product_15(498) <= '0';
partial_product_15(499) <= '0';
partial_product_15(500) <= '0';
partial_product_15(501) <= '0';
partial_product_15(502) <= '0';
partial_product_15(503) <= '0';
partial_product_15(504) <= '0';
partial_product_15(505) <= '0';
partial_product_15(506) <= '0';
partial_product_15(507) <= '0';
partial_product_15(508) <= '0';
partial_product_15(509) <= '0';
partial_product_15(510) <= '0';
partial_product_15(511) <= '0';
partial_product_15(512) <= '0';
partial_product_16(0) <= '0';
partial_product_16(1) <= '0';
partial_product_16(2) <= '0';
partial_product_16(3) <= '0';
partial_product_16(4) <= '0';
partial_product_16(5) <= '0';
partial_product_16(6) <= '0';
partial_product_16(7) <= '0';
partial_product_16(8) <= '0';
partial_product_16(9) <= '0';
partial_product_16(10) <= '0';
partial_product_16(11) <= '0';
partial_product_16(12) <= '0';
partial_product_16(13) <= '0';
partial_product_16(14) <= '0';
partial_product_16(15) <= '0';
partial_product_16(16) <= '0';
partial_product_16(17) <= '0';
partial_product_16(18) <= '0';
partial_product_16(19) <= '0';
partial_product_16(20) <= '0';
partial_product_16(21) <= '0';
partial_product_16(22) <= '0';
partial_product_16(23) <= '0';
partial_product_16(24) <= '0';
partial_product_16(25) <= '0';
partial_product_16(26) <= '0';
partial_product_16(27) <= '0';
partial_product_16(28) <= '0';
partial_product_16(29) <= '0';
partial_product_16(30) <= '0';
partial_product_16(31) <= '0';
partial_product_16(32) <= '0';
partial_product_16(33) <= '0';
partial_product_16(34) <= '0';
partial_product_16(35) <= '0';
partial_product_16(36) <= '0';
partial_product_16(37) <= '0';
partial_product_16(38) <= '0';
partial_product_16(39) <= '0';
partial_product_16(40) <= '0';
partial_product_16(41) <= '0';
partial_product_16(42) <= '0';
partial_product_16(43) <= '0';
partial_product_16(44) <= '0';
partial_product_16(45) <= '0';
partial_product_16(46) <= '0';
partial_product_16(47) <= '0';
partial_product_16(48) <= '0';
partial_product_16(49) <= '0';
partial_product_16(50) <= '0';
partial_product_16(51) <= '0';
partial_product_16(52) <= '0';
partial_product_16(53) <= '0';
partial_product_16(54) <= '0';
partial_product_16(55) <= '0';
partial_product_16(56) <= '0';
partial_product_16(57) <= '0';
partial_product_16(58) <= '0';
partial_product_16(59) <= '0';
partial_product_16(60) <= '0';
partial_product_16(61) <= '0';
partial_product_16(62) <= '0';
partial_product_16(63) <= '0';
partial_product_16(64) <= '0';
partial_product_16(65) <= '0';
partial_product_16(66) <= '0';
partial_product_16(67) <= '0';
partial_product_16(68) <= '0';
partial_product_16(69) <= '0';
partial_product_16(70) <= '0';
partial_product_16(71) <= '0';
partial_product_16(72) <= '0';
partial_product_16(73) <= '0';
partial_product_16(74) <= '0';
partial_product_16(75) <= '0';
partial_product_16(76) <= '0';
partial_product_16(77) <= '0';
partial_product_16(78) <= '0';
partial_product_16(79) <= '0';
partial_product_16(80) <= '0';
partial_product_16(81) <= '0';
partial_product_16(82) <= '0';
partial_product_16(83) <= '0';
partial_product_16(84) <= '0';
partial_product_16(85) <= '0';
partial_product_16(86) <= '0';
partial_product_16(87) <= '0';
partial_product_16(88) <= '0';
partial_product_16(89) <= '0';
partial_product_16(90) <= '0';
partial_product_16(91) <= '0';
partial_product_16(92) <= '0';
partial_product_16(93) <= '0';
partial_product_16(94) <= '0';
partial_product_16(95) <= '0';
partial_product_16(96) <= '0';
partial_product_16(97) <= '0';
partial_product_16(98) <= '0';
partial_product_16(99) <= '0';
partial_product_16(100) <= '0';
partial_product_16(101) <= '0';
partial_product_16(102) <= '0';
partial_product_16(103) <= '0';
partial_product_16(104) <= '0';
partial_product_16(105) <= '0';
partial_product_16(106) <= '0';
partial_product_16(107) <= '0';
partial_product_16(108) <= '0';
partial_product_16(109) <= '0';
partial_product_16(110) <= '0';
partial_product_16(111) <= '0';
partial_product_16(112) <= '0';
partial_product_16(113) <= '0';
partial_product_16(114) <= '0';
partial_product_16(115) <= '0';
partial_product_16(116) <= '0';
partial_product_16(117) <= '0';
partial_product_16(118) <= '0';
partial_product_16(119) <= '0';
partial_product_16(120) <= '0';
partial_product_16(121) <= '0';
partial_product_16(122) <= '0';
partial_product_16(123) <= '0';
partial_product_16(124) <= '0';
partial_product_16(125) <= '0';
partial_product_16(126) <= '0';
partial_product_16(127) <= '0';
partial_product_16(128) <= '0';
partial_product_16(129) <= '0';
partial_product_16(130) <= '0';
partial_product_16(131) <= '0';
partial_product_16(132) <= '0';
partial_product_16(133) <= '0';
partial_product_16(134) <= '0';
partial_product_16(135) <= '0';
partial_product_16(136) <= '0';
partial_product_16(137) <= '0';
partial_product_16(138) <= '0';
partial_product_16(139) <= '0';
partial_product_16(140) <= '0';
partial_product_16(141) <= '0';
partial_product_16(142) <= '0';
partial_product_16(143) <= '0';
partial_product_16(144) <= '0';
partial_product_16(145) <= '0';
partial_product_16(146) <= '0';
partial_product_16(147) <= '0';
partial_product_16(148) <= '0';
partial_product_16(149) <= '0';
partial_product_16(150) <= '0';
partial_product_16(151) <= '0';
partial_product_16(152) <= '0';
partial_product_16(153) <= '0';
partial_product_16(154) <= '0';
partial_product_16(155) <= '0';
partial_product_16(156) <= '0';
partial_product_16(157) <= '0';
partial_product_16(158) <= '0';
partial_product_16(159) <= '0';
partial_product_16(160) <= '0';
partial_product_16(161) <= '0';
partial_product_16(162) <= '0';
partial_product_16(163) <= '0';
partial_product_16(164) <= '0';
partial_product_16(165) <= '0';
partial_product_16(166) <= '0';
partial_product_16(167) <= '0';
partial_product_16(168) <= temp_mult_56(168);
partial_product_16(169) <= temp_mult_56(169);
partial_product_16(170) <= temp_mult_56(170);
partial_product_16(171) <= temp_mult_56(171);
partial_product_16(172) <= temp_mult_56(172);
partial_product_16(173) <= temp_mult_56(173);
partial_product_16(174) <= temp_mult_56(174);
partial_product_16(175) <= temp_mult_56(175);
partial_product_16(176) <= temp_mult_56(176);
partial_product_16(177) <= temp_mult_56(177);
partial_product_16(178) <= temp_mult_56(178);
partial_product_16(179) <= temp_mult_56(179);
partial_product_16(180) <= temp_mult_56(180);
partial_product_16(181) <= temp_mult_56(181);
partial_product_16(182) <= temp_mult_56(182);
partial_product_16(183) <= temp_mult_56(183);
partial_product_16(184) <= temp_mult_56(184);
partial_product_16(185) <= temp_mult_56(185);
partial_product_16(186) <= temp_mult_56(186);
partial_product_16(187) <= temp_mult_56(187);
partial_product_16(188) <= temp_mult_56(188);
partial_product_16(189) <= temp_mult_56(189);
partial_product_16(190) <= temp_mult_56(190);
partial_product_16(191) <= temp_mult_56(191);
partial_product_16(192) <= temp_mult_56(192);
partial_product_16(193) <= temp_mult_56(193);
partial_product_16(194) <= temp_mult_56(194);
partial_product_16(195) <= temp_mult_56(195);
partial_product_16(196) <= temp_mult_56(196);
partial_product_16(197) <= temp_mult_56(197);
partial_product_16(198) <= temp_mult_56(198);
partial_product_16(199) <= temp_mult_56(199);
partial_product_16(200) <= temp_mult_56(200);
partial_product_16(201) <= temp_mult_56(201);
partial_product_16(202) <= temp_mult_56(202);
partial_product_16(203) <= temp_mult_56(203);
partial_product_16(204) <= temp_mult_56(204);
partial_product_16(205) <= temp_mult_56(205);
partial_product_16(206) <= temp_mult_56(206);
partial_product_16(207) <= temp_mult_56(207);
partial_product_16(208) <= temp_mult_56(208);
partial_product_16(209) <= temp_mult_65(209);
partial_product_16(210) <= temp_mult_65(210);
partial_product_16(211) <= temp_mult_65(211);
partial_product_16(212) <= temp_mult_65(212);
partial_product_16(213) <= temp_mult_65(213);
partial_product_16(214) <= temp_mult_65(214);
partial_product_16(215) <= temp_mult_65(215);
partial_product_16(216) <= temp_mult_65(216);
partial_product_16(217) <= temp_mult_65(217);
partial_product_16(218) <= temp_mult_65(218);
partial_product_16(219) <= temp_mult_65(219);
partial_product_16(220) <= temp_mult_65(220);
partial_product_16(221) <= temp_mult_65(221);
partial_product_16(222) <= temp_mult_65(222);
partial_product_16(223) <= temp_mult_65(223);
partial_product_16(224) <= temp_mult_65(224);
partial_product_16(225) <= temp_mult_65(225);
partial_product_16(226) <= temp_mult_65(226);
partial_product_16(227) <= temp_mult_65(227);
partial_product_16(228) <= temp_mult_65(228);
partial_product_16(229) <= temp_mult_65(229);
partial_product_16(230) <= temp_mult_65(230);
partial_product_16(231) <= temp_mult_65(231);
partial_product_16(232) <= temp_mult_65(232);
partial_product_16(233) <= temp_mult_65(233);
partial_product_16(234) <= temp_mult_65(234);
partial_product_16(235) <= temp_mult_65(235);
partial_product_16(236) <= temp_mult_65(236);
partial_product_16(237) <= temp_mult_65(237);
partial_product_16(238) <= temp_mult_65(238);
partial_product_16(239) <= temp_mult_65(239);
partial_product_16(240) <= temp_mult_65(240);
partial_product_16(241) <= temp_mult_65(241);
partial_product_16(242) <= temp_mult_65(242);
partial_product_16(243) <= temp_mult_65(243);
partial_product_16(244) <= temp_mult_65(244);
partial_product_16(245) <= temp_mult_65(245);
partial_product_16(246) <= temp_mult_65(246);
partial_product_16(247) <= temp_mult_65(247);
partial_product_16(248) <= temp_mult_65(248);
partial_product_16(249) <= temp_mult_65(249);
partial_product_16(250) <= temp_mult_74(250);
partial_product_16(251) <= temp_mult_74(251);
partial_product_16(252) <= temp_mult_74(252);
partial_product_16(253) <= temp_mult_74(253);
partial_product_16(254) <= temp_mult_74(254);
partial_product_16(255) <= temp_mult_74(255);
partial_product_16(256) <= temp_mult_74(256);
partial_product_16(257) <= temp_mult_74(257);
partial_product_16(258) <= temp_mult_74(258);
partial_product_16(259) <= temp_mult_74(259);
partial_product_16(260) <= temp_mult_74(260);
partial_product_16(261) <= temp_mult_74(261);
partial_product_16(262) <= temp_mult_74(262);
partial_product_16(263) <= temp_mult_74(263);
partial_product_16(264) <= temp_mult_74(264);
partial_product_16(265) <= temp_mult_74(265);
partial_product_16(266) <= temp_mult_74(266);
partial_product_16(267) <= temp_mult_74(267);
partial_product_16(268) <= temp_mult_74(268);
partial_product_16(269) <= temp_mult_74(269);
partial_product_16(270) <= temp_mult_74(270);
partial_product_16(271) <= temp_mult_74(271);
partial_product_16(272) <= temp_mult_74(272);
partial_product_16(273) <= temp_mult_74(273);
partial_product_16(274) <= temp_mult_74(274);
partial_product_16(275) <= temp_mult_74(275);
partial_product_16(276) <= temp_mult_74(276);
partial_product_16(277) <= temp_mult_74(277);
partial_product_16(278) <= temp_mult_74(278);
partial_product_16(279) <= temp_mult_74(279);
partial_product_16(280) <= temp_mult_74(280);
partial_product_16(281) <= temp_mult_74(281);
partial_product_16(282) <= temp_mult_74(282);
partial_product_16(283) <= temp_mult_74(283);
partial_product_16(284) <= temp_mult_74(284);
partial_product_16(285) <= temp_mult_74(285);
partial_product_16(286) <= temp_mult_74(286);
partial_product_16(287) <= temp_mult_74(287);
partial_product_16(288) <= temp_mult_74(288);
partial_product_16(289) <= temp_mult_74(289);
partial_product_16(290) <= temp_mult_74(290);
partial_product_16(291) <= '0';
partial_product_16(292) <= '0';
partial_product_16(293) <= temp_mult_109(293);
partial_product_16(294) <= temp_mult_109(294);
partial_product_16(295) <= temp_mult_109(295);
partial_product_16(296) <= temp_mult_109(296);
partial_product_16(297) <= temp_mult_109(297);
partial_product_16(298) <= temp_mult_109(298);
partial_product_16(299) <= temp_mult_109(299);
partial_product_16(300) <= temp_mult_109(300);
partial_product_16(301) <= temp_mult_109(301);
partial_product_16(302) <= temp_mult_109(302);
partial_product_16(303) <= temp_mult_109(303);
partial_product_16(304) <= temp_mult_109(304);
partial_product_16(305) <= temp_mult_109(305);
partial_product_16(306) <= temp_mult_109(306);
partial_product_16(307) <= temp_mult_109(307);
partial_product_16(308) <= temp_mult_109(308);
partial_product_16(309) <= temp_mult_109(309);
partial_product_16(310) <= temp_mult_109(310);
partial_product_16(311) <= temp_mult_109(311);
partial_product_16(312) <= temp_mult_109(312);
partial_product_16(313) <= temp_mult_109(313);
partial_product_16(314) <= temp_mult_109(314);
partial_product_16(315) <= temp_mult_109(315);
partial_product_16(316) <= temp_mult_109(316);
partial_product_16(317) <= temp_mult_109(317);
partial_product_16(318) <= temp_mult_109(318);
partial_product_16(319) <= temp_mult_109(319);
partial_product_16(320) <= temp_mult_109(320);
partial_product_16(321) <= temp_mult_109(321);
partial_product_16(322) <= temp_mult_109(322);
partial_product_16(323) <= temp_mult_109(323);
partial_product_16(324) <= temp_mult_109(324);
partial_product_16(325) <= temp_mult_109(325);
partial_product_16(326) <= temp_mult_109(326);
partial_product_16(327) <= temp_mult_109(327);
partial_product_16(328) <= temp_mult_109(328);
partial_product_16(329) <= temp_mult_109(329);
partial_product_16(330) <= temp_mult_109(330);
partial_product_16(331) <= temp_mult_109(331);
partial_product_16(332) <= temp_mult_109(332);
partial_product_16(333) <= temp_mult_109(333);
partial_product_16(334) <= temp_mult_118(334);
partial_product_16(335) <= temp_mult_118(335);
partial_product_16(336) <= temp_mult_118(336);
partial_product_16(337) <= temp_mult_118(337);
partial_product_16(338) <= temp_mult_118(338);
partial_product_16(339) <= temp_mult_118(339);
partial_product_16(340) <= temp_mult_118(340);
partial_product_16(341) <= temp_mult_118(341);
partial_product_16(342) <= temp_mult_118(342);
partial_product_16(343) <= temp_mult_118(343);
partial_product_16(344) <= temp_mult_118(344);
partial_product_16(345) <= temp_mult_118(345);
partial_product_16(346) <= temp_mult_118(346);
partial_product_16(347) <= temp_mult_118(347);
partial_product_16(348) <= temp_mult_118(348);
partial_product_16(349) <= temp_mult_118(349);
partial_product_16(350) <= temp_mult_118(350);
partial_product_16(351) <= temp_mult_118(351);
partial_product_16(352) <= temp_mult_118(352);
partial_product_16(353) <= temp_mult_118(353);
partial_product_16(354) <= temp_mult_118(354);
partial_product_16(355) <= temp_mult_118(355);
partial_product_16(356) <= temp_mult_118(356);
partial_product_16(357) <= temp_mult_118(357);
partial_product_16(358) <= temp_mult_118(358);
partial_product_16(359) <= temp_mult_118(359);
partial_product_16(360) <= temp_mult_118(360);
partial_product_16(361) <= temp_mult_118(361);
partial_product_16(362) <= temp_mult_118(362);
partial_product_16(363) <= temp_mult_118(363);
partial_product_16(364) <= temp_mult_118(364);
partial_product_16(365) <= temp_mult_118(365);
partial_product_16(366) <= temp_mult_118(366);
partial_product_16(367) <= temp_mult_118(367);
partial_product_16(368) <= temp_mult_118(368);
partial_product_16(369) <= temp_mult_118(369);
partial_product_16(370) <= temp_mult_118(370);
partial_product_16(371) <= temp_mult_118(371);
partial_product_16(372) <= temp_mult_118(372);
partial_product_16(373) <= temp_mult_118(373);
partial_product_16(374) <= temp_mult_118(374);
partial_product_16(375) <= '0';
partial_product_16(376) <= '0';
partial_product_16(377) <= '0';
partial_product_16(378) <= '0';
partial_product_16(379) <= '0';
partial_product_16(380) <= '0';
partial_product_16(381) <= '0';
partial_product_16(382) <= '0';
partial_product_16(383) <= '0';
partial_product_16(384) <= '0';
partial_product_16(385) <= '0';
partial_product_16(386) <= '0';
partial_product_16(387) <= '0';
partial_product_16(388) <= '0';
partial_product_16(389) <= '0';
partial_product_16(390) <= '0';
partial_product_16(391) <= '0';
partial_product_16(392) <= '0';
partial_product_16(393) <= '0';
partial_product_16(394) <= '0';
partial_product_16(395) <= '0';
partial_product_16(396) <= '0';
partial_product_16(397) <= '0';
partial_product_16(398) <= '0';
partial_product_16(399) <= '0';
partial_product_16(400) <= '0';
partial_product_16(401) <= '0';
partial_product_16(402) <= '0';
partial_product_16(403) <= '0';
partial_product_16(404) <= '0';
partial_product_16(405) <= '0';
partial_product_16(406) <= '0';
partial_product_16(407) <= '0';
partial_product_16(408) <= '0';
partial_product_16(409) <= '0';
partial_product_16(410) <= '0';
partial_product_16(411) <= '0';
partial_product_16(412) <= '0';
partial_product_16(413) <= '0';
partial_product_16(414) <= '0';
partial_product_16(415) <= '0';
partial_product_16(416) <= '0';
partial_product_16(417) <= '0';
partial_product_16(418) <= '0';
partial_product_16(419) <= '0';
partial_product_16(420) <= '0';
partial_product_16(421) <= '0';
partial_product_16(422) <= '0';
partial_product_16(423) <= '0';
partial_product_16(424) <= '0';
partial_product_16(425) <= '0';
partial_product_16(426) <= '0';
partial_product_16(427) <= '0';
partial_product_16(428) <= '0';
partial_product_16(429) <= '0';
partial_product_16(430) <= '0';
partial_product_16(431) <= '0';
partial_product_16(432) <= '0';
partial_product_16(433) <= '0';
partial_product_16(434) <= '0';
partial_product_16(435) <= '0';
partial_product_16(436) <= '0';
partial_product_16(437) <= '0';
partial_product_16(438) <= '0';
partial_product_16(439) <= '0';
partial_product_16(440) <= '0';
partial_product_16(441) <= '0';
partial_product_16(442) <= '0';
partial_product_16(443) <= '0';
partial_product_16(444) <= '0';
partial_product_16(445) <= '0';
partial_product_16(446) <= '0';
partial_product_16(447) <= '0';
partial_product_16(448) <= '0';
partial_product_16(449) <= '0';
partial_product_16(450) <= '0';
partial_product_16(451) <= '0';
partial_product_16(452) <= '0';
partial_product_16(453) <= '0';
partial_product_16(454) <= '0';
partial_product_16(455) <= '0';
partial_product_16(456) <= '0';
partial_product_16(457) <= '0';
partial_product_16(458) <= '0';
partial_product_16(459) <= '0';
partial_product_16(460) <= '0';
partial_product_16(461) <= '0';
partial_product_16(462) <= '0';
partial_product_16(463) <= '0';
partial_product_16(464) <= '0';
partial_product_16(465) <= '0';
partial_product_16(466) <= '0';
partial_product_16(467) <= '0';
partial_product_16(468) <= '0';
partial_product_16(469) <= '0';
partial_product_16(470) <= '0';
partial_product_16(471) <= '0';
partial_product_16(472) <= '0';
partial_product_16(473) <= '0';
partial_product_16(474) <= '0';
partial_product_16(475) <= '0';
partial_product_16(476) <= '0';
partial_product_16(477) <= '0';
partial_product_16(478) <= '0';
partial_product_16(479) <= '0';
partial_product_16(480) <= '0';
partial_product_16(481) <= '0';
partial_product_16(482) <= '0';
partial_product_16(483) <= '0';
partial_product_16(484) <= '0';
partial_product_16(485) <= '0';
partial_product_16(486) <= '0';
partial_product_16(487) <= '0';
partial_product_16(488) <= '0';
partial_product_16(489) <= '0';
partial_product_16(490) <= '0';
partial_product_16(491) <= '0';
partial_product_16(492) <= '0';
partial_product_16(493) <= '0';
partial_product_16(494) <= '0';
partial_product_16(495) <= '0';
partial_product_16(496) <= '0';
partial_product_16(497) <= '0';
partial_product_16(498) <= '0';
partial_product_16(499) <= '0';
partial_product_16(500) <= '0';
partial_product_16(501) <= '0';
partial_product_16(502) <= '0';
partial_product_16(503) <= '0';
partial_product_16(504) <= '0';
partial_product_16(505) <= '0';
partial_product_16(506) <= '0';
partial_product_16(507) <= '0';
partial_product_16(508) <= '0';
partial_product_16(509) <= '0';
partial_product_16(510) <= '0';
partial_product_16(511) <= '0';
partial_product_16(512) <= '0';
partial_product_17(0) <= '0';
partial_product_17(1) <= '0';
partial_product_17(2) <= '0';
partial_product_17(3) <= '0';
partial_product_17(4) <= '0';
partial_product_17(5) <= '0';
partial_product_17(6) <= '0';
partial_product_17(7) <= '0';
partial_product_17(8) <= '0';
partial_product_17(9) <= '0';
partial_product_17(10) <= '0';
partial_product_17(11) <= '0';
partial_product_17(12) <= '0';
partial_product_17(13) <= '0';
partial_product_17(14) <= '0';
partial_product_17(15) <= '0';
partial_product_17(16) <= '0';
partial_product_17(17) <= '0';
partial_product_17(18) <= '0';
partial_product_17(19) <= '0';
partial_product_17(20) <= '0';
partial_product_17(21) <= '0';
partial_product_17(22) <= '0';
partial_product_17(23) <= '0';
partial_product_17(24) <= '0';
partial_product_17(25) <= '0';
partial_product_17(26) <= '0';
partial_product_17(27) <= '0';
partial_product_17(28) <= '0';
partial_product_17(29) <= '0';
partial_product_17(30) <= '0';
partial_product_17(31) <= '0';
partial_product_17(32) <= '0';
partial_product_17(33) <= '0';
partial_product_17(34) <= '0';
partial_product_17(35) <= '0';
partial_product_17(36) <= '0';
partial_product_17(37) <= '0';
partial_product_17(38) <= '0';
partial_product_17(39) <= '0';
partial_product_17(40) <= '0';
partial_product_17(41) <= '0';
partial_product_17(42) <= '0';
partial_product_17(43) <= '0';
partial_product_17(44) <= '0';
partial_product_17(45) <= '0';
partial_product_17(46) <= '0';
partial_product_17(47) <= '0';
partial_product_17(48) <= '0';
partial_product_17(49) <= '0';
partial_product_17(50) <= '0';
partial_product_17(51) <= '0';
partial_product_17(52) <= '0';
partial_product_17(53) <= '0';
partial_product_17(54) <= '0';
partial_product_17(55) <= '0';
partial_product_17(56) <= '0';
partial_product_17(57) <= '0';
partial_product_17(58) <= '0';
partial_product_17(59) <= '0';
partial_product_17(60) <= '0';
partial_product_17(61) <= '0';
partial_product_17(62) <= '0';
partial_product_17(63) <= '0';
partial_product_17(64) <= '0';
partial_product_17(65) <= '0';
partial_product_17(66) <= '0';
partial_product_17(67) <= '0';
partial_product_17(68) <= '0';
partial_product_17(69) <= '0';
partial_product_17(70) <= '0';
partial_product_17(71) <= '0';
partial_product_17(72) <= '0';
partial_product_17(73) <= '0';
partial_product_17(74) <= '0';
partial_product_17(75) <= '0';
partial_product_17(76) <= '0';
partial_product_17(77) <= '0';
partial_product_17(78) <= '0';
partial_product_17(79) <= '0';
partial_product_17(80) <= '0';
partial_product_17(81) <= '0';
partial_product_17(82) <= '0';
partial_product_17(83) <= '0';
partial_product_17(84) <= '0';
partial_product_17(85) <= '0';
partial_product_17(86) <= '0';
partial_product_17(87) <= '0';
partial_product_17(88) <= '0';
partial_product_17(89) <= '0';
partial_product_17(90) <= '0';
partial_product_17(91) <= '0';
partial_product_17(92) <= '0';
partial_product_17(93) <= '0';
partial_product_17(94) <= '0';
partial_product_17(95) <= '0';
partial_product_17(96) <= '0';
partial_product_17(97) <= '0';
partial_product_17(98) <= '0';
partial_product_17(99) <= '0';
partial_product_17(100) <= '0';
partial_product_17(101) <= '0';
partial_product_17(102) <= '0';
partial_product_17(103) <= '0';
partial_product_17(104) <= '0';
partial_product_17(105) <= '0';
partial_product_17(106) <= '0';
partial_product_17(107) <= '0';
partial_product_17(108) <= '0';
partial_product_17(109) <= '0';
partial_product_17(110) <= '0';
partial_product_17(111) <= '0';
partial_product_17(112) <= '0';
partial_product_17(113) <= '0';
partial_product_17(114) <= '0';
partial_product_17(115) <= '0';
partial_product_17(116) <= '0';
partial_product_17(117) <= '0';
partial_product_17(118) <= '0';
partial_product_17(119) <= '0';
partial_product_17(120) <= '0';
partial_product_17(121) <= '0';
partial_product_17(122) <= '0';
partial_product_17(123) <= '0';
partial_product_17(124) <= '0';
partial_product_17(125) <= '0';
partial_product_17(126) <= '0';
partial_product_17(127) <= '0';
partial_product_17(128) <= '0';
partial_product_17(129) <= '0';
partial_product_17(130) <= '0';
partial_product_17(131) <= '0';
partial_product_17(132) <= '0';
partial_product_17(133) <= '0';
partial_product_17(134) <= '0';
partial_product_17(135) <= '0';
partial_product_17(136) <= '0';
partial_product_17(137) <= '0';
partial_product_17(138) <= '0';
partial_product_17(139) <= '0';
partial_product_17(140) <= '0';
partial_product_17(141) <= '0';
partial_product_17(142) <= '0';
partial_product_17(143) <= '0';
partial_product_17(144) <= '0';
partial_product_17(145) <= '0';
partial_product_17(146) <= '0';
partial_product_17(147) <= '0';
partial_product_17(148) <= '0';
partial_product_17(149) <= '0';
partial_product_17(150) <= '0';
partial_product_17(151) <= '0';
partial_product_17(152) <= '0';
partial_product_17(153) <= '0';
partial_product_17(154) <= '0';
partial_product_17(155) <= '0';
partial_product_17(156) <= '0';
partial_product_17(157) <= '0';
partial_product_17(158) <= '0';
partial_product_17(159) <= '0';
partial_product_17(160) <= '0';
partial_product_17(161) <= '0';
partial_product_17(162) <= '0';
partial_product_17(163) <= '0';
partial_product_17(164) <= '0';
partial_product_17(165) <= '0';
partial_product_17(166) <= '0';
partial_product_17(167) <= '0';
partial_product_17(168) <= '0';
partial_product_17(169) <= '0';
partial_product_17(170) <= temp_mult_82(170);
partial_product_17(171) <= temp_mult_82(171);
partial_product_17(172) <= temp_mult_82(172);
partial_product_17(173) <= temp_mult_82(173);
partial_product_17(174) <= temp_mult_82(174);
partial_product_17(175) <= temp_mult_82(175);
partial_product_17(176) <= temp_mult_82(176);
partial_product_17(177) <= temp_mult_82(177);
partial_product_17(178) <= temp_mult_82(178);
partial_product_17(179) <= temp_mult_82(179);
partial_product_17(180) <= temp_mult_82(180);
partial_product_17(181) <= temp_mult_82(181);
partial_product_17(182) <= temp_mult_82(182);
partial_product_17(183) <= temp_mult_82(183);
partial_product_17(184) <= temp_mult_82(184);
partial_product_17(185) <= temp_mult_82(185);
partial_product_17(186) <= temp_mult_82(186);
partial_product_17(187) <= temp_mult_82(187);
partial_product_17(188) <= temp_mult_82(188);
partial_product_17(189) <= temp_mult_82(189);
partial_product_17(190) <= temp_mult_82(190);
partial_product_17(191) <= temp_mult_82(191);
partial_product_17(192) <= temp_mult_82(192);
partial_product_17(193) <= temp_mult_82(193);
partial_product_17(194) <= temp_mult_82(194);
partial_product_17(195) <= temp_mult_82(195);
partial_product_17(196) <= temp_mult_82(196);
partial_product_17(197) <= temp_mult_82(197);
partial_product_17(198) <= temp_mult_82(198);
partial_product_17(199) <= temp_mult_82(199);
partial_product_17(200) <= temp_mult_82(200);
partial_product_17(201) <= temp_mult_82(201);
partial_product_17(202) <= temp_mult_82(202);
partial_product_17(203) <= temp_mult_82(203);
partial_product_17(204) <= temp_mult_82(204);
partial_product_17(205) <= temp_mult_82(205);
partial_product_17(206) <= temp_mult_82(206);
partial_product_17(207) <= temp_mult_82(207);
partial_product_17(208) <= temp_mult_82(208);
partial_product_17(209) <= temp_mult_82(209);
partial_product_17(210) <= temp_mult_82(210);
partial_product_17(211) <= temp_mult_91(211);
partial_product_17(212) <= temp_mult_91(212);
partial_product_17(213) <= temp_mult_91(213);
partial_product_17(214) <= temp_mult_91(214);
partial_product_17(215) <= temp_mult_91(215);
partial_product_17(216) <= temp_mult_91(216);
partial_product_17(217) <= temp_mult_91(217);
partial_product_17(218) <= temp_mult_91(218);
partial_product_17(219) <= temp_mult_91(219);
partial_product_17(220) <= temp_mult_91(220);
partial_product_17(221) <= temp_mult_91(221);
partial_product_17(222) <= temp_mult_91(222);
partial_product_17(223) <= temp_mult_91(223);
partial_product_17(224) <= temp_mult_91(224);
partial_product_17(225) <= temp_mult_91(225);
partial_product_17(226) <= temp_mult_91(226);
partial_product_17(227) <= temp_mult_91(227);
partial_product_17(228) <= temp_mult_91(228);
partial_product_17(229) <= temp_mult_91(229);
partial_product_17(230) <= temp_mult_91(230);
partial_product_17(231) <= temp_mult_91(231);
partial_product_17(232) <= temp_mult_91(232);
partial_product_17(233) <= temp_mult_91(233);
partial_product_17(234) <= temp_mult_91(234);
partial_product_17(235) <= temp_mult_91(235);
partial_product_17(236) <= temp_mult_91(236);
partial_product_17(237) <= temp_mult_91(237);
partial_product_17(238) <= temp_mult_91(238);
partial_product_17(239) <= temp_mult_91(239);
partial_product_17(240) <= temp_mult_91(240);
partial_product_17(241) <= temp_mult_91(241);
partial_product_17(242) <= temp_mult_91(242);
partial_product_17(243) <= temp_mult_91(243);
partial_product_17(244) <= temp_mult_91(244);
partial_product_17(245) <= temp_mult_91(245);
partial_product_17(246) <= temp_mult_91(246);
partial_product_17(247) <= temp_mult_91(247);
partial_product_17(248) <= temp_mult_91(248);
partial_product_17(249) <= temp_mult_91(249);
partial_product_17(250) <= temp_mult_91(250);
partial_product_17(251) <= temp_mult_91(251);
partial_product_17(252) <= temp_mult_100(252);
partial_product_17(253) <= temp_mult_100(253);
partial_product_17(254) <= temp_mult_100(254);
partial_product_17(255) <= temp_mult_100(255);
partial_product_17(256) <= temp_mult_100(256);
partial_product_17(257) <= temp_mult_100(257);
partial_product_17(258) <= temp_mult_100(258);
partial_product_17(259) <= temp_mult_100(259);
partial_product_17(260) <= temp_mult_100(260);
partial_product_17(261) <= temp_mult_100(261);
partial_product_17(262) <= temp_mult_100(262);
partial_product_17(263) <= temp_mult_100(263);
partial_product_17(264) <= temp_mult_100(264);
partial_product_17(265) <= temp_mult_100(265);
partial_product_17(266) <= temp_mult_100(266);
partial_product_17(267) <= temp_mult_100(267);
partial_product_17(268) <= temp_mult_100(268);
partial_product_17(269) <= temp_mult_100(269);
partial_product_17(270) <= temp_mult_100(270);
partial_product_17(271) <= temp_mult_100(271);
partial_product_17(272) <= temp_mult_100(272);
partial_product_17(273) <= temp_mult_100(273);
partial_product_17(274) <= temp_mult_100(274);
partial_product_17(275) <= temp_mult_100(275);
partial_product_17(276) <= temp_mult_100(276);
partial_product_17(277) <= temp_mult_100(277);
partial_product_17(278) <= temp_mult_100(278);
partial_product_17(279) <= temp_mult_100(279);
partial_product_17(280) <= temp_mult_100(280);
partial_product_17(281) <= temp_mult_100(281);
partial_product_17(282) <= temp_mult_100(282);
partial_product_17(283) <= temp_mult_100(283);
partial_product_17(284) <= temp_mult_100(284);
partial_product_17(285) <= temp_mult_100(285);
partial_product_17(286) <= temp_mult_100(286);
partial_product_17(287) <= temp_mult_100(287);
partial_product_17(288) <= temp_mult_100(288);
partial_product_17(289) <= temp_mult_100(289);
partial_product_17(290) <= temp_mult_100(290);
partial_product_17(291) <= temp_mult_100(291);
partial_product_17(292) <= temp_mult_100(292);
partial_product_17(293) <= '0';
partial_product_17(294) <= '0';
partial_product_17(295) <= '0';
partial_product_17(296) <= '0';
partial_product_17(297) <= '0';
partial_product_17(298) <= '0';
partial_product_17(299) <= '0';
partial_product_17(300) <= '0';
partial_product_17(301) <= '0';
partial_product_17(302) <= '0';
partial_product_17(303) <= temp_mult_103(303);
partial_product_17(304) <= temp_mult_103(304);
partial_product_17(305) <= temp_mult_103(305);
partial_product_17(306) <= temp_mult_103(306);
partial_product_17(307) <= temp_mult_103(307);
partial_product_17(308) <= temp_mult_103(308);
partial_product_17(309) <= temp_mult_103(309);
partial_product_17(310) <= temp_mult_103(310);
partial_product_17(311) <= temp_mult_103(311);
partial_product_17(312) <= temp_mult_103(312);
partial_product_17(313) <= temp_mult_103(313);
partial_product_17(314) <= temp_mult_103(314);
partial_product_17(315) <= temp_mult_103(315);
partial_product_17(316) <= temp_mult_103(316);
partial_product_17(317) <= temp_mult_103(317);
partial_product_17(318) <= temp_mult_103(318);
partial_product_17(319) <= temp_mult_103(319);
partial_product_17(320) <= temp_mult_103(320);
partial_product_17(321) <= temp_mult_103(321);
partial_product_17(322) <= temp_mult_103(322);
partial_product_17(323) <= temp_mult_103(323);
partial_product_17(324) <= temp_mult_103(324);
partial_product_17(325) <= temp_mult_103(325);
partial_product_17(326) <= temp_mult_103(326);
partial_product_17(327) <= temp_mult_103(327);
partial_product_17(328) <= temp_mult_103(328);
partial_product_17(329) <= temp_mult_103(329);
partial_product_17(330) <= temp_mult_103(330);
partial_product_17(331) <= temp_mult_103(331);
partial_product_17(332) <= temp_mult_103(332);
partial_product_17(333) <= temp_mult_103(333);
partial_product_17(334) <= temp_mult_103(334);
partial_product_17(335) <= temp_mult_103(335);
partial_product_17(336) <= temp_mult_103(336);
partial_product_17(337) <= temp_mult_103(337);
partial_product_17(338) <= temp_mult_103(338);
partial_product_17(339) <= temp_mult_103(339);
partial_product_17(340) <= temp_mult_103(340);
partial_product_17(341) <= temp_mult_103(341);
partial_product_17(342) <= temp_mult_103(342);
partial_product_17(343) <= temp_mult_103(343);
partial_product_17(344) <= '0';
partial_product_17(345) <= '0';
partial_product_17(346) <= '0';
partial_product_17(347) <= '0';
partial_product_17(348) <= '0';
partial_product_17(349) <= '0';
partial_product_17(350) <= '0';
partial_product_17(351) <= '0';
partial_product_17(352) <= '0';
partial_product_17(353) <= '0';
partial_product_17(354) <= '0';
partial_product_17(355) <= '0';
partial_product_17(356) <= '0';
partial_product_17(357) <= '0';
partial_product_17(358) <= '0';
partial_product_17(359) <= '0';
partial_product_17(360) <= '0';
partial_product_17(361) <= '0';
partial_product_17(362) <= '0';
partial_product_17(363) <= '0';
partial_product_17(364) <= '0';
partial_product_17(365) <= '0';
partial_product_17(366) <= '0';
partial_product_17(367) <= '0';
partial_product_17(368) <= '0';
partial_product_17(369) <= '0';
partial_product_17(370) <= '0';
partial_product_17(371) <= '0';
partial_product_17(372) <= '0';
partial_product_17(373) <= '0';
partial_product_17(374) <= '0';
partial_product_17(375) <= '0';
partial_product_17(376) <= '0';
partial_product_17(377) <= '0';
partial_product_17(378) <= '0';
partial_product_17(379) <= '0';
partial_product_17(380) <= '0';
partial_product_17(381) <= '0';
partial_product_17(382) <= '0';
partial_product_17(383) <= '0';
partial_product_17(384) <= '0';
partial_product_17(385) <= '0';
partial_product_17(386) <= '0';
partial_product_17(387) <= '0';
partial_product_17(388) <= '0';
partial_product_17(389) <= '0';
partial_product_17(390) <= '0';
partial_product_17(391) <= '0';
partial_product_17(392) <= '0';
partial_product_17(393) <= '0';
partial_product_17(394) <= '0';
partial_product_17(395) <= '0';
partial_product_17(396) <= '0';
partial_product_17(397) <= '0';
partial_product_17(398) <= '0';
partial_product_17(399) <= '0';
partial_product_17(400) <= '0';
partial_product_17(401) <= '0';
partial_product_17(402) <= '0';
partial_product_17(403) <= '0';
partial_product_17(404) <= '0';
partial_product_17(405) <= '0';
partial_product_17(406) <= '0';
partial_product_17(407) <= '0';
partial_product_17(408) <= '0';
partial_product_17(409) <= '0';
partial_product_17(410) <= '0';
partial_product_17(411) <= '0';
partial_product_17(412) <= '0';
partial_product_17(413) <= '0';
partial_product_17(414) <= '0';
partial_product_17(415) <= '0';
partial_product_17(416) <= '0';
partial_product_17(417) <= '0';
partial_product_17(418) <= '0';
partial_product_17(419) <= '0';
partial_product_17(420) <= '0';
partial_product_17(421) <= '0';
partial_product_17(422) <= '0';
partial_product_17(423) <= '0';
partial_product_17(424) <= '0';
partial_product_17(425) <= '0';
partial_product_17(426) <= '0';
partial_product_17(427) <= '0';
partial_product_17(428) <= '0';
partial_product_17(429) <= '0';
partial_product_17(430) <= '0';
partial_product_17(431) <= '0';
partial_product_17(432) <= '0';
partial_product_17(433) <= '0';
partial_product_17(434) <= '0';
partial_product_17(435) <= '0';
partial_product_17(436) <= '0';
partial_product_17(437) <= '0';
partial_product_17(438) <= '0';
partial_product_17(439) <= '0';
partial_product_17(440) <= '0';
partial_product_17(441) <= '0';
partial_product_17(442) <= '0';
partial_product_17(443) <= '0';
partial_product_17(444) <= '0';
partial_product_17(445) <= '0';
partial_product_17(446) <= '0';
partial_product_17(447) <= '0';
partial_product_17(448) <= '0';
partial_product_17(449) <= '0';
partial_product_17(450) <= '0';
partial_product_17(451) <= '0';
partial_product_17(452) <= '0';
partial_product_17(453) <= '0';
partial_product_17(454) <= '0';
partial_product_17(455) <= '0';
partial_product_17(456) <= '0';
partial_product_17(457) <= '0';
partial_product_17(458) <= '0';
partial_product_17(459) <= '0';
partial_product_17(460) <= '0';
partial_product_17(461) <= '0';
partial_product_17(462) <= '0';
partial_product_17(463) <= '0';
partial_product_17(464) <= '0';
partial_product_17(465) <= '0';
partial_product_17(466) <= '0';
partial_product_17(467) <= '0';
partial_product_17(468) <= '0';
partial_product_17(469) <= '0';
partial_product_17(470) <= '0';
partial_product_17(471) <= '0';
partial_product_17(472) <= '0';
partial_product_17(473) <= '0';
partial_product_17(474) <= '0';
partial_product_17(475) <= '0';
partial_product_17(476) <= '0';
partial_product_17(477) <= '0';
partial_product_17(478) <= '0';
partial_product_17(479) <= '0';
partial_product_17(480) <= '0';
partial_product_17(481) <= '0';
partial_product_17(482) <= '0';
partial_product_17(483) <= '0';
partial_product_17(484) <= '0';
partial_product_17(485) <= '0';
partial_product_17(486) <= '0';
partial_product_17(487) <= '0';
partial_product_17(488) <= '0';
partial_product_17(489) <= '0';
partial_product_17(490) <= '0';
partial_product_17(491) <= '0';
partial_product_17(492) <= '0';
partial_product_17(493) <= '0';
partial_product_17(494) <= '0';
partial_product_17(495) <= '0';
partial_product_17(496) <= '0';
partial_product_17(497) <= '0';
partial_product_17(498) <= '0';
partial_product_17(499) <= '0';
partial_product_17(500) <= '0';
partial_product_17(501) <= '0';
partial_product_17(502) <= '0';
partial_product_17(503) <= '0';
partial_product_17(504) <= '0';
partial_product_17(505) <= '0';
partial_product_17(506) <= '0';
partial_product_17(507) <= '0';
partial_product_17(508) <= '0';
partial_product_17(509) <= '0';
partial_product_17(510) <= '0';
partial_product_17(511) <= '0';
partial_product_17(512) <= '0';
partial_product_18(0) <= '0';
partial_product_18(1) <= '0';
partial_product_18(2) <= '0';
partial_product_18(3) <= '0';
partial_product_18(4) <= '0';
partial_product_18(5) <= '0';
partial_product_18(6) <= '0';
partial_product_18(7) <= '0';
partial_product_18(8) <= '0';
partial_product_18(9) <= '0';
partial_product_18(10) <= '0';
partial_product_18(11) <= '0';
partial_product_18(12) <= '0';
partial_product_18(13) <= '0';
partial_product_18(14) <= '0';
partial_product_18(15) <= '0';
partial_product_18(16) <= '0';
partial_product_18(17) <= '0';
partial_product_18(18) <= '0';
partial_product_18(19) <= '0';
partial_product_18(20) <= '0';
partial_product_18(21) <= '0';
partial_product_18(22) <= '0';
partial_product_18(23) <= '0';
partial_product_18(24) <= '0';
partial_product_18(25) <= '0';
partial_product_18(26) <= '0';
partial_product_18(27) <= '0';
partial_product_18(28) <= '0';
partial_product_18(29) <= '0';
partial_product_18(30) <= '0';
partial_product_18(31) <= '0';
partial_product_18(32) <= '0';
partial_product_18(33) <= '0';
partial_product_18(34) <= '0';
partial_product_18(35) <= '0';
partial_product_18(36) <= '0';
partial_product_18(37) <= '0';
partial_product_18(38) <= '0';
partial_product_18(39) <= '0';
partial_product_18(40) <= '0';
partial_product_18(41) <= '0';
partial_product_18(42) <= '0';
partial_product_18(43) <= '0';
partial_product_18(44) <= '0';
partial_product_18(45) <= '0';
partial_product_18(46) <= '0';
partial_product_18(47) <= '0';
partial_product_18(48) <= '0';
partial_product_18(49) <= '0';
partial_product_18(50) <= '0';
partial_product_18(51) <= '0';
partial_product_18(52) <= '0';
partial_product_18(53) <= '0';
partial_product_18(54) <= '0';
partial_product_18(55) <= '0';
partial_product_18(56) <= '0';
partial_product_18(57) <= '0';
partial_product_18(58) <= '0';
partial_product_18(59) <= '0';
partial_product_18(60) <= '0';
partial_product_18(61) <= '0';
partial_product_18(62) <= '0';
partial_product_18(63) <= '0';
partial_product_18(64) <= '0';
partial_product_18(65) <= '0';
partial_product_18(66) <= '0';
partial_product_18(67) <= '0';
partial_product_18(68) <= '0';
partial_product_18(69) <= '0';
partial_product_18(70) <= '0';
partial_product_18(71) <= '0';
partial_product_18(72) <= '0';
partial_product_18(73) <= '0';
partial_product_18(74) <= '0';
partial_product_18(75) <= '0';
partial_product_18(76) <= '0';
partial_product_18(77) <= '0';
partial_product_18(78) <= '0';
partial_product_18(79) <= '0';
partial_product_18(80) <= '0';
partial_product_18(81) <= '0';
partial_product_18(82) <= '0';
partial_product_18(83) <= '0';
partial_product_18(84) <= '0';
partial_product_18(85) <= '0';
partial_product_18(86) <= '0';
partial_product_18(87) <= '0';
partial_product_18(88) <= '0';
partial_product_18(89) <= '0';
partial_product_18(90) <= '0';
partial_product_18(91) <= '0';
partial_product_18(92) <= '0';
partial_product_18(93) <= '0';
partial_product_18(94) <= '0';
partial_product_18(95) <= '0';
partial_product_18(96) <= '0';
partial_product_18(97) <= '0';
partial_product_18(98) <= '0';
partial_product_18(99) <= '0';
partial_product_18(100) <= '0';
partial_product_18(101) <= '0';
partial_product_18(102) <= '0';
partial_product_18(103) <= '0';
partial_product_18(104) <= '0';
partial_product_18(105) <= '0';
partial_product_18(106) <= '0';
partial_product_18(107) <= '0';
partial_product_18(108) <= '0';
partial_product_18(109) <= '0';
partial_product_18(110) <= '0';
partial_product_18(111) <= '0';
partial_product_18(112) <= '0';
partial_product_18(113) <= '0';
partial_product_18(114) <= '0';
partial_product_18(115) <= '0';
partial_product_18(116) <= '0';
partial_product_18(117) <= '0';
partial_product_18(118) <= '0';
partial_product_18(119) <= '0';
partial_product_18(120) <= '0';
partial_product_18(121) <= '0';
partial_product_18(122) <= '0';
partial_product_18(123) <= '0';
partial_product_18(124) <= '0';
partial_product_18(125) <= '0';
partial_product_18(126) <= '0';
partial_product_18(127) <= '0';
partial_product_18(128) <= '0';
partial_product_18(129) <= '0';
partial_product_18(130) <= '0';
partial_product_18(131) <= '0';
partial_product_18(132) <= '0';
partial_product_18(133) <= '0';
partial_product_18(134) <= '0';
partial_product_18(135) <= '0';
partial_product_18(136) <= '0';
partial_product_18(137) <= '0';
partial_product_18(138) <= '0';
partial_product_18(139) <= '0';
partial_product_18(140) <= '0';
partial_product_18(141) <= '0';
partial_product_18(142) <= '0';
partial_product_18(143) <= '0';
partial_product_18(144) <= '0';
partial_product_18(145) <= '0';
partial_product_18(146) <= '0';
partial_product_18(147) <= '0';
partial_product_18(148) <= '0';
partial_product_18(149) <= '0';
partial_product_18(150) <= '0';
partial_product_18(151) <= '0';
partial_product_18(152) <= '0';
partial_product_18(153) <= '0';
partial_product_18(154) <= '0';
partial_product_18(155) <= '0';
partial_product_18(156) <= '0';
partial_product_18(157) <= '0';
partial_product_18(158) <= '0';
partial_product_18(159) <= '0';
partial_product_18(160) <= '0';
partial_product_18(161) <= '0';
partial_product_18(162) <= '0';
partial_product_18(163) <= '0';
partial_product_18(164) <= '0';
partial_product_18(165) <= '0';
partial_product_18(166) <= '0';
partial_product_18(167) <= '0';
partial_product_18(168) <= '0';
partial_product_18(169) <= '0';
partial_product_18(170) <= '0';
partial_product_18(171) <= '0';
partial_product_18(172) <= '0';
partial_product_18(173) <= '0';
partial_product_18(174) <= '0';
partial_product_18(175) <= '0';
partial_product_18(176) <= '0';
partial_product_18(177) <= '0';
partial_product_18(178) <= '0';
partial_product_18(179) <= '0';
partial_product_18(180) <= '0';
partial_product_18(181) <= '0';
partial_product_18(182) <= '0';
partial_product_18(183) <= '0';
partial_product_18(184) <= '0';
partial_product_18(185) <= '0';
partial_product_18(186) <= '0';
partial_product_18(187) <= temp_mult_83(187);
partial_product_18(188) <= temp_mult_83(188);
partial_product_18(189) <= temp_mult_83(189);
partial_product_18(190) <= temp_mult_83(190);
partial_product_18(191) <= temp_mult_83(191);
partial_product_18(192) <= temp_mult_83(192);
partial_product_18(193) <= temp_mult_83(193);
partial_product_18(194) <= temp_mult_83(194);
partial_product_18(195) <= temp_mult_83(195);
partial_product_18(196) <= temp_mult_83(196);
partial_product_18(197) <= temp_mult_83(197);
partial_product_18(198) <= temp_mult_83(198);
partial_product_18(199) <= temp_mult_83(199);
partial_product_18(200) <= temp_mult_83(200);
partial_product_18(201) <= temp_mult_83(201);
partial_product_18(202) <= temp_mult_83(202);
partial_product_18(203) <= temp_mult_83(203);
partial_product_18(204) <= temp_mult_83(204);
partial_product_18(205) <= temp_mult_83(205);
partial_product_18(206) <= temp_mult_83(206);
partial_product_18(207) <= temp_mult_83(207);
partial_product_18(208) <= temp_mult_83(208);
partial_product_18(209) <= temp_mult_83(209);
partial_product_18(210) <= temp_mult_83(210);
partial_product_18(211) <= temp_mult_83(211);
partial_product_18(212) <= temp_mult_83(212);
partial_product_18(213) <= temp_mult_83(213);
partial_product_18(214) <= temp_mult_83(214);
partial_product_18(215) <= temp_mult_83(215);
partial_product_18(216) <= temp_mult_83(216);
partial_product_18(217) <= temp_mult_83(217);
partial_product_18(218) <= temp_mult_83(218);
partial_product_18(219) <= temp_mult_83(219);
partial_product_18(220) <= temp_mult_83(220);
partial_product_18(221) <= temp_mult_83(221);
partial_product_18(222) <= temp_mult_83(222);
partial_product_18(223) <= temp_mult_83(223);
partial_product_18(224) <= temp_mult_83(224);
partial_product_18(225) <= temp_mult_83(225);
partial_product_18(226) <= temp_mult_83(226);
partial_product_18(227) <= temp_mult_83(227);
partial_product_18(228) <= temp_mult_92(228);
partial_product_18(229) <= temp_mult_92(229);
partial_product_18(230) <= temp_mult_92(230);
partial_product_18(231) <= temp_mult_92(231);
partial_product_18(232) <= temp_mult_92(232);
partial_product_18(233) <= temp_mult_92(233);
partial_product_18(234) <= temp_mult_92(234);
partial_product_18(235) <= temp_mult_92(235);
partial_product_18(236) <= temp_mult_92(236);
partial_product_18(237) <= temp_mult_92(237);
partial_product_18(238) <= temp_mult_92(238);
partial_product_18(239) <= temp_mult_92(239);
partial_product_18(240) <= temp_mult_92(240);
partial_product_18(241) <= temp_mult_92(241);
partial_product_18(242) <= temp_mult_92(242);
partial_product_18(243) <= temp_mult_92(243);
partial_product_18(244) <= temp_mult_92(244);
partial_product_18(245) <= temp_mult_92(245);
partial_product_18(246) <= temp_mult_92(246);
partial_product_18(247) <= temp_mult_92(247);
partial_product_18(248) <= temp_mult_92(248);
partial_product_18(249) <= temp_mult_92(249);
partial_product_18(250) <= temp_mult_92(250);
partial_product_18(251) <= temp_mult_92(251);
partial_product_18(252) <= temp_mult_92(252);
partial_product_18(253) <= temp_mult_92(253);
partial_product_18(254) <= temp_mult_92(254);
partial_product_18(255) <= temp_mult_92(255);
partial_product_18(256) <= temp_mult_92(256);
partial_product_18(257) <= temp_mult_92(257);
partial_product_18(258) <= temp_mult_92(258);
partial_product_18(259) <= temp_mult_92(259);
partial_product_18(260) <= temp_mult_92(260);
partial_product_18(261) <= temp_mult_92(261);
partial_product_18(262) <= temp_mult_92(262);
partial_product_18(263) <= temp_mult_92(263);
partial_product_18(264) <= temp_mult_92(264);
partial_product_18(265) <= temp_mult_92(265);
partial_product_18(266) <= temp_mult_92(266);
partial_product_18(267) <= temp_mult_92(267);
partial_product_18(268) <= temp_mult_92(268);
partial_product_18(269) <= temp_mult_101(269);
partial_product_18(270) <= temp_mult_101(270);
partial_product_18(271) <= temp_mult_101(271);
partial_product_18(272) <= temp_mult_101(272);
partial_product_18(273) <= temp_mult_101(273);
partial_product_18(274) <= temp_mult_101(274);
partial_product_18(275) <= temp_mult_101(275);
partial_product_18(276) <= temp_mult_101(276);
partial_product_18(277) <= temp_mult_101(277);
partial_product_18(278) <= temp_mult_101(278);
partial_product_18(279) <= temp_mult_101(279);
partial_product_18(280) <= temp_mult_101(280);
partial_product_18(281) <= temp_mult_101(281);
partial_product_18(282) <= temp_mult_101(282);
partial_product_18(283) <= temp_mult_101(283);
partial_product_18(284) <= temp_mult_101(284);
partial_product_18(285) <= temp_mult_101(285);
partial_product_18(286) <= temp_mult_101(286);
partial_product_18(287) <= temp_mult_101(287);
partial_product_18(288) <= temp_mult_101(288);
partial_product_18(289) <= temp_mult_101(289);
partial_product_18(290) <= temp_mult_101(290);
partial_product_18(291) <= temp_mult_101(291);
partial_product_18(292) <= temp_mult_101(292);
partial_product_18(293) <= temp_mult_101(293);
partial_product_18(294) <= temp_mult_101(294);
partial_product_18(295) <= temp_mult_101(295);
partial_product_18(296) <= temp_mult_101(296);
partial_product_18(297) <= temp_mult_101(297);
partial_product_18(298) <= temp_mult_101(298);
partial_product_18(299) <= temp_mult_101(299);
partial_product_18(300) <= temp_mult_101(300);
partial_product_18(301) <= temp_mult_101(301);
partial_product_18(302) <= temp_mult_101(302);
partial_product_18(303) <= temp_mult_101(303);
partial_product_18(304) <= temp_mult_101(304);
partial_product_18(305) <= temp_mult_101(305);
partial_product_18(306) <= temp_mult_101(306);
partial_product_18(307) <= temp_mult_101(307);
partial_product_18(308) <= temp_mult_101(308);
partial_product_18(309) <= temp_mult_101(309);
partial_product_18(310) <= '0';
partial_product_18(311) <= '0';
partial_product_18(312) <= '0';
partial_product_18(313) <= '0';
partial_product_18(314) <= '0';
partial_product_18(315) <= '0';
partial_product_18(316) <= '0';
partial_product_18(317) <= '0';
partial_product_18(318) <= '0';
partial_product_18(319) <= '0';
partial_product_18(320) <= '0';
partial_product_18(321) <= '0';
partial_product_18(322) <= '0';
partial_product_18(323) <= '0';
partial_product_18(324) <= '0';
partial_product_18(325) <= '0';
partial_product_18(326) <= '0';
partial_product_18(327) <= '0';
partial_product_18(328) <= '0';
partial_product_18(329) <= '0';
partial_product_18(330) <= '0';
partial_product_18(331) <= '0';
partial_product_18(332) <= '0';
partial_product_18(333) <= '0';
partial_product_18(334) <= '0';
partial_product_18(335) <= '0';
partial_product_18(336) <= '0';
partial_product_18(337) <= '0';
partial_product_18(338) <= '0';
partial_product_18(339) <= '0';
partial_product_18(340) <= '0';
partial_product_18(341) <= '0';
partial_product_18(342) <= '0';
partial_product_18(343) <= '0';
partial_product_18(344) <= '0';
partial_product_18(345) <= '0';
partial_product_18(346) <= '0';
partial_product_18(347) <= '0';
partial_product_18(348) <= '0';
partial_product_18(349) <= '0';
partial_product_18(350) <= '0';
partial_product_18(351) <= '0';
partial_product_18(352) <= '0';
partial_product_18(353) <= '0';
partial_product_18(354) <= '0';
partial_product_18(355) <= '0';
partial_product_18(356) <= '0';
partial_product_18(357) <= '0';
partial_product_18(358) <= '0';
partial_product_18(359) <= '0';
partial_product_18(360) <= '0';
partial_product_18(361) <= '0';
partial_product_18(362) <= '0';
partial_product_18(363) <= '0';
partial_product_18(364) <= '0';
partial_product_18(365) <= '0';
partial_product_18(366) <= '0';
partial_product_18(367) <= '0';
partial_product_18(368) <= '0';
partial_product_18(369) <= '0';
partial_product_18(370) <= '0';
partial_product_18(371) <= '0';
partial_product_18(372) <= '0';
partial_product_18(373) <= '0';
partial_product_18(374) <= '0';
partial_product_18(375) <= '0';
partial_product_18(376) <= '0';
partial_product_18(377) <= '0';
partial_product_18(378) <= '0';
partial_product_18(379) <= '0';
partial_product_18(380) <= '0';
partial_product_18(381) <= '0';
partial_product_18(382) <= '0';
partial_product_18(383) <= '0';
partial_product_18(384) <= '0';
partial_product_18(385) <= '0';
partial_product_18(386) <= '0';
partial_product_18(387) <= '0';
partial_product_18(388) <= '0';
partial_product_18(389) <= '0';
partial_product_18(390) <= '0';
partial_product_18(391) <= '0';
partial_product_18(392) <= '0';
partial_product_18(393) <= '0';
partial_product_18(394) <= '0';
partial_product_18(395) <= '0';
partial_product_18(396) <= '0';
partial_product_18(397) <= '0';
partial_product_18(398) <= '0';
partial_product_18(399) <= '0';
partial_product_18(400) <= '0';
partial_product_18(401) <= '0';
partial_product_18(402) <= '0';
partial_product_18(403) <= '0';
partial_product_18(404) <= '0';
partial_product_18(405) <= '0';
partial_product_18(406) <= '0';
partial_product_18(407) <= '0';
partial_product_18(408) <= '0';
partial_product_18(409) <= '0';
partial_product_18(410) <= '0';
partial_product_18(411) <= '0';
partial_product_18(412) <= '0';
partial_product_18(413) <= '0';
partial_product_18(414) <= '0';
partial_product_18(415) <= '0';
partial_product_18(416) <= '0';
partial_product_18(417) <= '0';
partial_product_18(418) <= '0';
partial_product_18(419) <= '0';
partial_product_18(420) <= '0';
partial_product_18(421) <= '0';
partial_product_18(422) <= '0';
partial_product_18(423) <= '0';
partial_product_18(424) <= '0';
partial_product_18(425) <= '0';
partial_product_18(426) <= '0';
partial_product_18(427) <= '0';
partial_product_18(428) <= '0';
partial_product_18(429) <= '0';
partial_product_18(430) <= '0';
partial_product_18(431) <= '0';
partial_product_18(432) <= '0';
partial_product_18(433) <= '0';
partial_product_18(434) <= '0';
partial_product_18(435) <= '0';
partial_product_18(436) <= '0';
partial_product_18(437) <= '0';
partial_product_18(438) <= '0';
partial_product_18(439) <= '0';
partial_product_18(440) <= '0';
partial_product_18(441) <= '0';
partial_product_18(442) <= '0';
partial_product_18(443) <= '0';
partial_product_18(444) <= '0';
partial_product_18(445) <= '0';
partial_product_18(446) <= '0';
partial_product_18(447) <= '0';
partial_product_18(448) <= '0';
partial_product_18(449) <= '0';
partial_product_18(450) <= '0';
partial_product_18(451) <= '0';
partial_product_18(452) <= '0';
partial_product_18(453) <= '0';
partial_product_18(454) <= '0';
partial_product_18(455) <= '0';
partial_product_18(456) <= '0';
partial_product_18(457) <= '0';
partial_product_18(458) <= '0';
partial_product_18(459) <= '0';
partial_product_18(460) <= '0';
partial_product_18(461) <= '0';
partial_product_18(462) <= '0';
partial_product_18(463) <= '0';
partial_product_18(464) <= '0';
partial_product_18(465) <= '0';
partial_product_18(466) <= '0';
partial_product_18(467) <= '0';
partial_product_18(468) <= '0';
partial_product_18(469) <= '0';
partial_product_18(470) <= '0';
partial_product_18(471) <= '0';
partial_product_18(472) <= '0';
partial_product_18(473) <= '0';
partial_product_18(474) <= '0';
partial_product_18(475) <= '0';
partial_product_18(476) <= '0';
partial_product_18(477) <= '0';
partial_product_18(478) <= '0';
partial_product_18(479) <= '0';
partial_product_18(480) <= '0';
partial_product_18(481) <= '0';
partial_product_18(482) <= '0';
partial_product_18(483) <= '0';
partial_product_18(484) <= '0';
partial_product_18(485) <= '0';
partial_product_18(486) <= '0';
partial_product_18(487) <= '0';
partial_product_18(488) <= '0';
partial_product_18(489) <= '0';
partial_product_18(490) <= '0';
partial_product_18(491) <= '0';
partial_product_18(492) <= '0';
partial_product_18(493) <= '0';
partial_product_18(494) <= '0';
partial_product_18(495) <= '0';
partial_product_18(496) <= '0';
partial_product_18(497) <= '0';
partial_product_18(498) <= '0';
partial_product_18(499) <= '0';
partial_product_18(500) <= '0';
partial_product_18(501) <= '0';
partial_product_18(502) <= '0';
partial_product_18(503) <= '0';
partial_product_18(504) <= '0';
partial_product_18(505) <= '0';
partial_product_18(506) <= '0';
partial_product_18(507) <= '0';
partial_product_18(508) <= '0';
partial_product_18(509) <= '0';
partial_product_18(510) <= '0';
partial_product_18(511) <= '0';
partial_product_18(512) <= '0';
partial_product_19(0) <= '0';
partial_product_19(1) <= '0';
partial_product_19(2) <= '0';
partial_product_19(3) <= '0';
partial_product_19(4) <= '0';
partial_product_19(5) <= '0';
partial_product_19(6) <= '0';
partial_product_19(7) <= '0';
partial_product_19(8) <= '0';
partial_product_19(9) <= '0';
partial_product_19(10) <= '0';
partial_product_19(11) <= '0';
partial_product_19(12) <= '0';
partial_product_19(13) <= '0';
partial_product_19(14) <= '0';
partial_product_19(15) <= '0';
partial_product_19(16) <= '0';
partial_product_19(17) <= '0';
partial_product_19(18) <= '0';
partial_product_19(19) <= '0';
partial_product_19(20) <= '0';
partial_product_19(21) <= '0';
partial_product_19(22) <= '0';
partial_product_19(23) <= '0';
partial_product_19(24) <= '0';
partial_product_19(25) <= '0';
partial_product_19(26) <= '0';
partial_product_19(27) <= '0';
partial_product_19(28) <= '0';
partial_product_19(29) <= '0';
partial_product_19(30) <= '0';
partial_product_19(31) <= '0';
partial_product_19(32) <= '0';
partial_product_19(33) <= '0';
partial_product_19(34) <= '0';
partial_product_19(35) <= '0';
partial_product_19(36) <= '0';
partial_product_19(37) <= '0';
partial_product_19(38) <= '0';
partial_product_19(39) <= '0';
partial_product_19(40) <= '0';
partial_product_19(41) <= '0';
partial_product_19(42) <= '0';
partial_product_19(43) <= '0';
partial_product_19(44) <= '0';
partial_product_19(45) <= '0';
partial_product_19(46) <= '0';
partial_product_19(47) <= '0';
partial_product_19(48) <= '0';
partial_product_19(49) <= '0';
partial_product_19(50) <= '0';
partial_product_19(51) <= '0';
partial_product_19(52) <= '0';
partial_product_19(53) <= '0';
partial_product_19(54) <= '0';
partial_product_19(55) <= '0';
partial_product_19(56) <= '0';
partial_product_19(57) <= '0';
partial_product_19(58) <= '0';
partial_product_19(59) <= '0';
partial_product_19(60) <= '0';
partial_product_19(61) <= '0';
partial_product_19(62) <= '0';
partial_product_19(63) <= '0';
partial_product_19(64) <= '0';
partial_product_19(65) <= '0';
partial_product_19(66) <= '0';
partial_product_19(67) <= '0';
partial_product_19(68) <= '0';
partial_product_19(69) <= '0';
partial_product_19(70) <= '0';
partial_product_19(71) <= '0';
partial_product_19(72) <= '0';
partial_product_19(73) <= '0';
partial_product_19(74) <= '0';
partial_product_19(75) <= '0';
partial_product_19(76) <= '0';
partial_product_19(77) <= '0';
partial_product_19(78) <= '0';
partial_product_19(79) <= '0';
partial_product_19(80) <= '0';
partial_product_19(81) <= '0';
partial_product_19(82) <= '0';
partial_product_19(83) <= '0';
partial_product_19(84) <= '0';
partial_product_19(85) <= '0';
partial_product_19(86) <= '0';
partial_product_19(87) <= '0';
partial_product_19(88) <= '0';
partial_product_19(89) <= '0';
partial_product_19(90) <= '0';
partial_product_19(91) <= '0';
partial_product_19(92) <= '0';
partial_product_19(93) <= '0';
partial_product_19(94) <= '0';
partial_product_19(95) <= '0';
partial_product_19(96) <= '0';
partial_product_19(97) <= '0';
partial_product_19(98) <= '0';
partial_product_19(99) <= '0';
partial_product_19(100) <= '0';
partial_product_19(101) <= '0';
partial_product_19(102) <= '0';
partial_product_19(103) <= '0';
partial_product_19(104) <= '0';
partial_product_19(105) <= '0';
partial_product_19(106) <= '0';
partial_product_19(107) <= '0';
partial_product_19(108) <= '0';
partial_product_19(109) <= '0';
partial_product_19(110) <= '0';
partial_product_19(111) <= '0';
partial_product_19(112) <= '0';
partial_product_19(113) <= '0';
partial_product_19(114) <= '0';
partial_product_19(115) <= '0';
partial_product_19(116) <= '0';
partial_product_19(117) <= '0';
partial_product_19(118) <= '0';
partial_product_19(119) <= '0';
partial_product_19(120) <= '0';
partial_product_19(121) <= '0';
partial_product_19(122) <= '0';
partial_product_19(123) <= '0';
partial_product_19(124) <= '0';
partial_product_19(125) <= '0';
partial_product_19(126) <= '0';
partial_product_19(127) <= '0';
partial_product_19(128) <= '0';
partial_product_19(129) <= '0';
partial_product_19(130) <= '0';
partial_product_19(131) <= '0';
partial_product_19(132) <= '0';
partial_product_19(133) <= '0';
partial_product_19(134) <= '0';
partial_product_19(135) <= '0';
partial_product_19(136) <= '0';
partial_product_19(137) <= '0';
partial_product_19(138) <= '0';
partial_product_19(139) <= '0';
partial_product_19(140) <= '0';
partial_product_19(141) <= '0';
partial_product_19(142) <= '0';
partial_product_19(143) <= '0';
partial_product_19(144) <= '0';
partial_product_19(145) <= '0';
partial_product_19(146) <= '0';
partial_product_19(147) <= '0';
partial_product_19(148) <= '0';
partial_product_19(149) <= '0';
partial_product_19(150) <= '0';
partial_product_19(151) <= '0';
partial_product_19(152) <= '0';
partial_product_19(153) <= '0';
partial_product_19(154) <= '0';
partial_product_19(155) <= '0';
partial_product_19(156) <= '0';
partial_product_19(157) <= '0';
partial_product_19(158) <= '0';
partial_product_19(159) <= '0';
partial_product_19(160) <= '0';
partial_product_19(161) <= '0';
partial_product_19(162) <= '0';
partial_product_19(163) <= '0';
partial_product_19(164) <= '0';
partial_product_19(165) <= '0';
partial_product_19(166) <= '0';
partial_product_19(167) <= '0';
partial_product_19(168) <= '0';
partial_product_19(169) <= '0';
partial_product_19(170) <= '0';
partial_product_19(171) <= '0';
partial_product_19(172) <= '0';
partial_product_19(173) <= '0';
partial_product_19(174) <= '0';
partial_product_19(175) <= '0';
partial_product_19(176) <= '0';
partial_product_19(177) <= '0';
partial_product_19(178) <= '0';
partial_product_19(179) <= '0';
partial_product_19(180) <= '0';
partial_product_19(181) <= '0';
partial_product_19(182) <= '0';
partial_product_19(183) <= '0';
partial_product_19(184) <= '0';
partial_product_19(185) <= '0';
partial_product_19(186) <= '0';
partial_product_19(187) <= '0';
partial_product_19(188) <= '0';
partial_product_19(189) <= '0';
partial_product_19(190) <= '0';
partial_product_19(191) <= '0';
partial_product_19(192) <= temp_mult_64(192);
partial_product_19(193) <= temp_mult_64(193);
partial_product_19(194) <= temp_mult_64(194);
partial_product_19(195) <= temp_mult_64(195);
partial_product_19(196) <= temp_mult_64(196);
partial_product_19(197) <= temp_mult_64(197);
partial_product_19(198) <= temp_mult_64(198);
partial_product_19(199) <= temp_mult_64(199);
partial_product_19(200) <= temp_mult_64(200);
partial_product_19(201) <= temp_mult_64(201);
partial_product_19(202) <= temp_mult_64(202);
partial_product_19(203) <= temp_mult_64(203);
partial_product_19(204) <= temp_mult_64(204);
partial_product_19(205) <= temp_mult_64(205);
partial_product_19(206) <= temp_mult_64(206);
partial_product_19(207) <= temp_mult_64(207);
partial_product_19(208) <= temp_mult_64(208);
partial_product_19(209) <= temp_mult_64(209);
partial_product_19(210) <= temp_mult_64(210);
partial_product_19(211) <= temp_mult_64(211);
partial_product_19(212) <= temp_mult_64(212);
partial_product_19(213) <= temp_mult_64(213);
partial_product_19(214) <= temp_mult_64(214);
partial_product_19(215) <= temp_mult_64(215);
partial_product_19(216) <= temp_mult_64(216);
partial_product_19(217) <= temp_mult_64(217);
partial_product_19(218) <= temp_mult_64(218);
partial_product_19(219) <= temp_mult_64(219);
partial_product_19(220) <= temp_mult_64(220);
partial_product_19(221) <= temp_mult_64(221);
partial_product_19(222) <= temp_mult_64(222);
partial_product_19(223) <= temp_mult_64(223);
partial_product_19(224) <= temp_mult_64(224);
partial_product_19(225) <= temp_mult_64(225);
partial_product_19(226) <= temp_mult_64(226);
partial_product_19(227) <= temp_mult_64(227);
partial_product_19(228) <= temp_mult_64(228);
partial_product_19(229) <= temp_mult_64(229);
partial_product_19(230) <= temp_mult_64(230);
partial_product_19(231) <= temp_mult_64(231);
partial_product_19(232) <= temp_mult_64(232);
partial_product_19(233) <= temp_mult_73(233);
partial_product_19(234) <= temp_mult_73(234);
partial_product_19(235) <= temp_mult_73(235);
partial_product_19(236) <= temp_mult_73(236);
partial_product_19(237) <= temp_mult_73(237);
partial_product_19(238) <= temp_mult_73(238);
partial_product_19(239) <= temp_mult_73(239);
partial_product_19(240) <= temp_mult_73(240);
partial_product_19(241) <= temp_mult_73(241);
partial_product_19(242) <= temp_mult_73(242);
partial_product_19(243) <= temp_mult_73(243);
partial_product_19(244) <= temp_mult_73(244);
partial_product_19(245) <= temp_mult_73(245);
partial_product_19(246) <= temp_mult_73(246);
partial_product_19(247) <= temp_mult_73(247);
partial_product_19(248) <= temp_mult_73(248);
partial_product_19(249) <= temp_mult_73(249);
partial_product_19(250) <= temp_mult_73(250);
partial_product_19(251) <= temp_mult_73(251);
partial_product_19(252) <= temp_mult_73(252);
partial_product_19(253) <= temp_mult_73(253);
partial_product_19(254) <= temp_mult_73(254);
partial_product_19(255) <= temp_mult_73(255);
partial_product_19(256) <= temp_mult_73(256);
partial_product_19(257) <= temp_mult_73(257);
partial_product_19(258) <= temp_mult_73(258);
partial_product_19(259) <= temp_mult_73(259);
partial_product_19(260) <= temp_mult_73(260);
partial_product_19(261) <= temp_mult_73(261);
partial_product_19(262) <= temp_mult_73(262);
partial_product_19(263) <= temp_mult_73(263);
partial_product_19(264) <= temp_mult_73(264);
partial_product_19(265) <= temp_mult_73(265);
partial_product_19(266) <= temp_mult_73(266);
partial_product_19(267) <= temp_mult_73(267);
partial_product_19(268) <= temp_mult_73(268);
partial_product_19(269) <= temp_mult_73(269);
partial_product_19(270) <= temp_mult_73(270);
partial_product_19(271) <= temp_mult_73(271);
partial_product_19(272) <= temp_mult_73(272);
partial_product_19(273) <= temp_mult_73(273);
partial_product_19(274) <= '0';
partial_product_19(275) <= '0';
partial_product_19(276) <= '0';
partial_product_19(277) <= '0';
partial_product_19(278) <= '0';
partial_product_19(279) <= temp_mult_95(279);
partial_product_19(280) <= temp_mult_95(280);
partial_product_19(281) <= temp_mult_95(281);
partial_product_19(282) <= temp_mult_95(282);
partial_product_19(283) <= temp_mult_95(283);
partial_product_19(284) <= temp_mult_95(284);
partial_product_19(285) <= temp_mult_95(285);
partial_product_19(286) <= temp_mult_95(286);
partial_product_19(287) <= temp_mult_95(287);
partial_product_19(288) <= temp_mult_95(288);
partial_product_19(289) <= temp_mult_95(289);
partial_product_19(290) <= temp_mult_95(290);
partial_product_19(291) <= temp_mult_95(291);
partial_product_19(292) <= temp_mult_95(292);
partial_product_19(293) <= temp_mult_95(293);
partial_product_19(294) <= temp_mult_95(294);
partial_product_19(295) <= temp_mult_95(295);
partial_product_19(296) <= temp_mult_95(296);
partial_product_19(297) <= temp_mult_95(297);
partial_product_19(298) <= temp_mult_95(298);
partial_product_19(299) <= temp_mult_95(299);
partial_product_19(300) <= temp_mult_95(300);
partial_product_19(301) <= temp_mult_95(301);
partial_product_19(302) <= temp_mult_95(302);
partial_product_19(303) <= temp_mult_95(303);
partial_product_19(304) <= temp_mult_95(304);
partial_product_19(305) <= temp_mult_95(305);
partial_product_19(306) <= temp_mult_95(306);
partial_product_19(307) <= temp_mult_95(307);
partial_product_19(308) <= temp_mult_95(308);
partial_product_19(309) <= temp_mult_95(309);
partial_product_19(310) <= temp_mult_95(310);
partial_product_19(311) <= temp_mult_95(311);
partial_product_19(312) <= temp_mult_95(312);
partial_product_19(313) <= temp_mult_95(313);
partial_product_19(314) <= temp_mult_95(314);
partial_product_19(315) <= temp_mult_95(315);
partial_product_19(316) <= temp_mult_95(316);
partial_product_19(317) <= temp_mult_95(317);
partial_product_19(318) <= temp_mult_95(318);
partial_product_19(319) <= temp_mult_95(319);
partial_product_19(320) <= '0';
partial_product_19(321) <= '0';
partial_product_19(322) <= '0';
partial_product_19(323) <= '0';
partial_product_19(324) <= '0';
partial_product_19(325) <= '0';
partial_product_19(326) <= '0';
partial_product_19(327) <= '0';
partial_product_19(328) <= '0';
partial_product_19(329) <= '0';
partial_product_19(330) <= '0';
partial_product_19(331) <= '0';
partial_product_19(332) <= '0';
partial_product_19(333) <= '0';
partial_product_19(334) <= '0';
partial_product_19(335) <= '0';
partial_product_19(336) <= '0';
partial_product_19(337) <= '0';
partial_product_19(338) <= '0';
partial_product_19(339) <= '0';
partial_product_19(340) <= '0';
partial_product_19(341) <= '0';
partial_product_19(342) <= '0';
partial_product_19(343) <= '0';
partial_product_19(344) <= '0';
partial_product_19(345) <= '0';
partial_product_19(346) <= '0';
partial_product_19(347) <= '0';
partial_product_19(348) <= '0';
partial_product_19(349) <= '0';
partial_product_19(350) <= '0';
partial_product_19(351) <= '0';
partial_product_19(352) <= '0';
partial_product_19(353) <= '0';
partial_product_19(354) <= '0';
partial_product_19(355) <= '0';
partial_product_19(356) <= '0';
partial_product_19(357) <= '0';
partial_product_19(358) <= '0';
partial_product_19(359) <= '0';
partial_product_19(360) <= '0';
partial_product_19(361) <= '0';
partial_product_19(362) <= '0';
partial_product_19(363) <= '0';
partial_product_19(364) <= '0';
partial_product_19(365) <= '0';
partial_product_19(366) <= '0';
partial_product_19(367) <= '0';
partial_product_19(368) <= '0';
partial_product_19(369) <= '0';
partial_product_19(370) <= '0';
partial_product_19(371) <= '0';
partial_product_19(372) <= '0';
partial_product_19(373) <= '0';
partial_product_19(374) <= '0';
partial_product_19(375) <= '0';
partial_product_19(376) <= '0';
partial_product_19(377) <= '0';
partial_product_19(378) <= '0';
partial_product_19(379) <= '0';
partial_product_19(380) <= '0';
partial_product_19(381) <= '0';
partial_product_19(382) <= '0';
partial_product_19(383) <= '0';
partial_product_19(384) <= '0';
partial_product_19(385) <= '0';
partial_product_19(386) <= '0';
partial_product_19(387) <= '0';
partial_product_19(388) <= '0';
partial_product_19(389) <= '0';
partial_product_19(390) <= '0';
partial_product_19(391) <= '0';
partial_product_19(392) <= '0';
partial_product_19(393) <= '0';
partial_product_19(394) <= '0';
partial_product_19(395) <= '0';
partial_product_19(396) <= '0';
partial_product_19(397) <= '0';
partial_product_19(398) <= '0';
partial_product_19(399) <= '0';
partial_product_19(400) <= '0';
partial_product_19(401) <= '0';
partial_product_19(402) <= '0';
partial_product_19(403) <= '0';
partial_product_19(404) <= '0';
partial_product_19(405) <= '0';
partial_product_19(406) <= '0';
partial_product_19(407) <= '0';
partial_product_19(408) <= '0';
partial_product_19(409) <= '0';
partial_product_19(410) <= '0';
partial_product_19(411) <= '0';
partial_product_19(412) <= '0';
partial_product_19(413) <= '0';
partial_product_19(414) <= '0';
partial_product_19(415) <= '0';
partial_product_19(416) <= '0';
partial_product_19(417) <= '0';
partial_product_19(418) <= '0';
partial_product_19(419) <= '0';
partial_product_19(420) <= '0';
partial_product_19(421) <= '0';
partial_product_19(422) <= '0';
partial_product_19(423) <= '0';
partial_product_19(424) <= '0';
partial_product_19(425) <= '0';
partial_product_19(426) <= '0';
partial_product_19(427) <= '0';
partial_product_19(428) <= '0';
partial_product_19(429) <= '0';
partial_product_19(430) <= '0';
partial_product_19(431) <= '0';
partial_product_19(432) <= '0';
partial_product_19(433) <= '0';
partial_product_19(434) <= '0';
partial_product_19(435) <= '0';
partial_product_19(436) <= '0';
partial_product_19(437) <= '0';
partial_product_19(438) <= '0';
partial_product_19(439) <= '0';
partial_product_19(440) <= '0';
partial_product_19(441) <= '0';
partial_product_19(442) <= '0';
partial_product_19(443) <= '0';
partial_product_19(444) <= '0';
partial_product_19(445) <= '0';
partial_product_19(446) <= '0';
partial_product_19(447) <= '0';
partial_product_19(448) <= '0';
partial_product_19(449) <= '0';
partial_product_19(450) <= '0';
partial_product_19(451) <= '0';
partial_product_19(452) <= '0';
partial_product_19(453) <= '0';
partial_product_19(454) <= '0';
partial_product_19(455) <= '0';
partial_product_19(456) <= '0';
partial_product_19(457) <= '0';
partial_product_19(458) <= '0';
partial_product_19(459) <= '0';
partial_product_19(460) <= '0';
partial_product_19(461) <= '0';
partial_product_19(462) <= '0';
partial_product_19(463) <= '0';
partial_product_19(464) <= '0';
partial_product_19(465) <= '0';
partial_product_19(466) <= '0';
partial_product_19(467) <= '0';
partial_product_19(468) <= '0';
partial_product_19(469) <= '0';
partial_product_19(470) <= '0';
partial_product_19(471) <= '0';
partial_product_19(472) <= '0';
partial_product_19(473) <= '0';
partial_product_19(474) <= '0';
partial_product_19(475) <= '0';
partial_product_19(476) <= '0';
partial_product_19(477) <= '0';
partial_product_19(478) <= '0';
partial_product_19(479) <= '0';
partial_product_19(480) <= '0';
partial_product_19(481) <= '0';
partial_product_19(482) <= '0';
partial_product_19(483) <= '0';
partial_product_19(484) <= '0';
partial_product_19(485) <= '0';
partial_product_19(486) <= '0';
partial_product_19(487) <= '0';
partial_product_19(488) <= '0';
partial_product_19(489) <= '0';
partial_product_19(490) <= '0';
partial_product_19(491) <= '0';
partial_product_19(492) <= '0';
partial_product_19(493) <= '0';
partial_product_19(494) <= '0';
partial_product_19(495) <= '0';
partial_product_19(496) <= '0';
partial_product_19(497) <= '0';
partial_product_19(498) <= '0';
partial_product_19(499) <= '0';
partial_product_19(500) <= '0';
partial_product_19(501) <= '0';
partial_product_19(502) <= '0';
partial_product_19(503) <= '0';
partial_product_19(504) <= '0';
partial_product_19(505) <= '0';
partial_product_19(506) <= '0';
partial_product_19(507) <= '0';
partial_product_19(508) <= '0';
partial_product_19(509) <= '0';
partial_product_19(510) <= '0';
partial_product_19(511) <= '0';
partial_product_19(512) <= '0';
partial_product_20(0) <= '0';
partial_product_20(1) <= '0';
partial_product_20(2) <= '0';
partial_product_20(3) <= '0';
partial_product_20(4) <= '0';
partial_product_20(5) <= '0';
partial_product_20(6) <= '0';
partial_product_20(7) <= '0';
partial_product_20(8) <= '0';
partial_product_20(9) <= '0';
partial_product_20(10) <= '0';
partial_product_20(11) <= '0';
partial_product_20(12) <= '0';
partial_product_20(13) <= '0';
partial_product_20(14) <= '0';
partial_product_20(15) <= '0';
partial_product_20(16) <= '0';
partial_product_20(17) <= '0';
partial_product_20(18) <= '0';
partial_product_20(19) <= '0';
partial_product_20(20) <= '0';
partial_product_20(21) <= '0';
partial_product_20(22) <= '0';
partial_product_20(23) <= '0';
partial_product_20(24) <= '0';
partial_product_20(25) <= '0';
partial_product_20(26) <= '0';
partial_product_20(27) <= '0';
partial_product_20(28) <= '0';
partial_product_20(29) <= '0';
partial_product_20(30) <= '0';
partial_product_20(31) <= '0';
partial_product_20(32) <= '0';
partial_product_20(33) <= '0';
partial_product_20(34) <= '0';
partial_product_20(35) <= '0';
partial_product_20(36) <= '0';
partial_product_20(37) <= '0';
partial_product_20(38) <= '0';
partial_product_20(39) <= '0';
partial_product_20(40) <= '0';
partial_product_20(41) <= '0';
partial_product_20(42) <= '0';
partial_product_20(43) <= '0';
partial_product_20(44) <= '0';
partial_product_20(45) <= '0';
partial_product_20(46) <= '0';
partial_product_20(47) <= '0';
partial_product_20(48) <= '0';
partial_product_20(49) <= '0';
partial_product_20(50) <= '0';
partial_product_20(51) <= '0';
partial_product_20(52) <= '0';
partial_product_20(53) <= '0';
partial_product_20(54) <= '0';
partial_product_20(55) <= '0';
partial_product_20(56) <= '0';
partial_product_20(57) <= '0';
partial_product_20(58) <= '0';
partial_product_20(59) <= '0';
partial_product_20(60) <= '0';
partial_product_20(61) <= '0';
partial_product_20(62) <= '0';
partial_product_20(63) <= '0';
partial_product_20(64) <= '0';
partial_product_20(65) <= '0';
partial_product_20(66) <= '0';
partial_product_20(67) <= '0';
partial_product_20(68) <= '0';
partial_product_20(69) <= '0';
partial_product_20(70) <= '0';
partial_product_20(71) <= '0';
partial_product_20(72) <= '0';
partial_product_20(73) <= '0';
partial_product_20(74) <= '0';
partial_product_20(75) <= '0';
partial_product_20(76) <= '0';
partial_product_20(77) <= '0';
partial_product_20(78) <= '0';
partial_product_20(79) <= '0';
partial_product_20(80) <= '0';
partial_product_20(81) <= '0';
partial_product_20(82) <= '0';
partial_product_20(83) <= '0';
partial_product_20(84) <= '0';
partial_product_20(85) <= '0';
partial_product_20(86) <= '0';
partial_product_20(87) <= '0';
partial_product_20(88) <= '0';
partial_product_20(89) <= '0';
partial_product_20(90) <= '0';
partial_product_20(91) <= '0';
partial_product_20(92) <= '0';
partial_product_20(93) <= '0';
partial_product_20(94) <= '0';
partial_product_20(95) <= '0';
partial_product_20(96) <= '0';
partial_product_20(97) <= '0';
partial_product_20(98) <= '0';
partial_product_20(99) <= '0';
partial_product_20(100) <= '0';
partial_product_20(101) <= '0';
partial_product_20(102) <= '0';
partial_product_20(103) <= '0';
partial_product_20(104) <= '0';
partial_product_20(105) <= '0';
partial_product_20(106) <= '0';
partial_product_20(107) <= '0';
partial_product_20(108) <= '0';
partial_product_20(109) <= '0';
partial_product_20(110) <= '0';
partial_product_20(111) <= '0';
partial_product_20(112) <= '0';
partial_product_20(113) <= '0';
partial_product_20(114) <= '0';
partial_product_20(115) <= '0';
partial_product_20(116) <= '0';
partial_product_20(117) <= '0';
partial_product_20(118) <= '0';
partial_product_20(119) <= '0';
partial_product_20(120) <= '0';
partial_product_20(121) <= '0';
partial_product_20(122) <= '0';
partial_product_20(123) <= '0';
partial_product_20(124) <= '0';
partial_product_20(125) <= '0';
partial_product_20(126) <= '0';
partial_product_20(127) <= '0';
partial_product_20(128) <= '0';
partial_product_20(129) <= '0';
partial_product_20(130) <= '0';
partial_product_20(131) <= '0';
partial_product_20(132) <= '0';
partial_product_20(133) <= '0';
partial_product_20(134) <= '0';
partial_product_20(135) <= '0';
partial_product_20(136) <= '0';
partial_product_20(137) <= '0';
partial_product_20(138) <= '0';
partial_product_20(139) <= '0';
partial_product_20(140) <= '0';
partial_product_20(141) <= '0';
partial_product_20(142) <= '0';
partial_product_20(143) <= '0';
partial_product_20(144) <= '0';
partial_product_20(145) <= '0';
partial_product_20(146) <= '0';
partial_product_20(147) <= '0';
partial_product_20(148) <= '0';
partial_product_20(149) <= '0';
partial_product_20(150) <= '0';
partial_product_20(151) <= '0';
partial_product_20(152) <= '0';
partial_product_20(153) <= '0';
partial_product_20(154) <= '0';
partial_product_20(155) <= '0';
partial_product_20(156) <= '0';
partial_product_20(157) <= '0';
partial_product_20(158) <= '0';
partial_product_20(159) <= '0';
partial_product_20(160) <= '0';
partial_product_20(161) <= '0';
partial_product_20(162) <= '0';
partial_product_20(163) <= '0';
partial_product_20(164) <= '0';
partial_product_20(165) <= '0';
partial_product_20(166) <= '0';
partial_product_20(167) <= '0';
partial_product_20(168) <= '0';
partial_product_20(169) <= '0';
partial_product_20(170) <= '0';
partial_product_20(171) <= '0';
partial_product_20(172) <= '0';
partial_product_20(173) <= '0';
partial_product_20(174) <= '0';
partial_product_20(175) <= '0';
partial_product_20(176) <= '0';
partial_product_20(177) <= '0';
partial_product_20(178) <= '0';
partial_product_20(179) <= '0';
partial_product_20(180) <= '0';
partial_product_20(181) <= '0';
partial_product_20(182) <= '0';
partial_product_20(183) <= '0';
partial_product_20(184) <= '0';
partial_product_20(185) <= '0';
partial_product_20(186) <= '0';
partial_product_20(187) <= '0';
partial_product_20(188) <= '0';
partial_product_20(189) <= '0';
partial_product_20(190) <= '0';
partial_product_20(191) <= '0';
partial_product_20(192) <= '0';
partial_product_20(193) <= '0';
partial_product_20(194) <= '0';
partial_product_20(195) <= '0';
partial_product_20(196) <= '0';
partial_product_20(197) <= '0';
partial_product_20(198) <= '0';
partial_product_20(199) <= '0';
partial_product_20(200) <= '0';
partial_product_20(201) <= '0';
partial_product_20(202) <= '0';
partial_product_20(203) <= '0';
partial_product_20(204) <= temp_mult_84(204);
partial_product_20(205) <= temp_mult_84(205);
partial_product_20(206) <= temp_mult_84(206);
partial_product_20(207) <= temp_mult_84(207);
partial_product_20(208) <= temp_mult_84(208);
partial_product_20(209) <= temp_mult_84(209);
partial_product_20(210) <= temp_mult_84(210);
partial_product_20(211) <= temp_mult_84(211);
partial_product_20(212) <= temp_mult_84(212);
partial_product_20(213) <= temp_mult_84(213);
partial_product_20(214) <= temp_mult_84(214);
partial_product_20(215) <= temp_mult_84(215);
partial_product_20(216) <= temp_mult_84(216);
partial_product_20(217) <= temp_mult_84(217);
partial_product_20(218) <= temp_mult_84(218);
partial_product_20(219) <= temp_mult_84(219);
partial_product_20(220) <= temp_mult_84(220);
partial_product_20(221) <= temp_mult_84(221);
partial_product_20(222) <= temp_mult_84(222);
partial_product_20(223) <= temp_mult_84(223);
partial_product_20(224) <= temp_mult_84(224);
partial_product_20(225) <= temp_mult_84(225);
partial_product_20(226) <= temp_mult_84(226);
partial_product_20(227) <= temp_mult_84(227);
partial_product_20(228) <= temp_mult_84(228);
partial_product_20(229) <= temp_mult_84(229);
partial_product_20(230) <= temp_mult_84(230);
partial_product_20(231) <= temp_mult_84(231);
partial_product_20(232) <= temp_mult_84(232);
partial_product_20(233) <= temp_mult_84(233);
partial_product_20(234) <= temp_mult_84(234);
partial_product_20(235) <= temp_mult_84(235);
partial_product_20(236) <= temp_mult_84(236);
partial_product_20(237) <= temp_mult_84(237);
partial_product_20(238) <= temp_mult_84(238);
partial_product_20(239) <= temp_mult_84(239);
partial_product_20(240) <= temp_mult_84(240);
partial_product_20(241) <= temp_mult_84(241);
partial_product_20(242) <= temp_mult_84(242);
partial_product_20(243) <= temp_mult_84(243);
partial_product_20(244) <= temp_mult_84(244);
partial_product_20(245) <= temp_mult_93(245);
partial_product_20(246) <= temp_mult_93(246);
partial_product_20(247) <= temp_mult_93(247);
partial_product_20(248) <= temp_mult_93(248);
partial_product_20(249) <= temp_mult_93(249);
partial_product_20(250) <= temp_mult_93(250);
partial_product_20(251) <= temp_mult_93(251);
partial_product_20(252) <= temp_mult_93(252);
partial_product_20(253) <= temp_mult_93(253);
partial_product_20(254) <= temp_mult_93(254);
partial_product_20(255) <= temp_mult_93(255);
partial_product_20(256) <= temp_mult_93(256);
partial_product_20(257) <= temp_mult_93(257);
partial_product_20(258) <= temp_mult_93(258);
partial_product_20(259) <= temp_mult_93(259);
partial_product_20(260) <= temp_mult_93(260);
partial_product_20(261) <= temp_mult_93(261);
partial_product_20(262) <= temp_mult_93(262);
partial_product_20(263) <= temp_mult_93(263);
partial_product_20(264) <= temp_mult_93(264);
partial_product_20(265) <= temp_mult_93(265);
partial_product_20(266) <= temp_mult_93(266);
partial_product_20(267) <= temp_mult_93(267);
partial_product_20(268) <= temp_mult_93(268);
partial_product_20(269) <= temp_mult_93(269);
partial_product_20(270) <= temp_mult_93(270);
partial_product_20(271) <= temp_mult_93(271);
partial_product_20(272) <= temp_mult_93(272);
partial_product_20(273) <= temp_mult_93(273);
partial_product_20(274) <= temp_mult_93(274);
partial_product_20(275) <= temp_mult_93(275);
partial_product_20(276) <= temp_mult_93(276);
partial_product_20(277) <= temp_mult_93(277);
partial_product_20(278) <= temp_mult_93(278);
partial_product_20(279) <= temp_mult_93(279);
partial_product_20(280) <= temp_mult_93(280);
partial_product_20(281) <= temp_mult_93(281);
partial_product_20(282) <= temp_mult_93(282);
partial_product_20(283) <= temp_mult_93(283);
partial_product_20(284) <= temp_mult_93(284);
partial_product_20(285) <= temp_mult_93(285);
partial_product_20(286) <= temp_mult_102(286);
partial_product_20(287) <= temp_mult_102(287);
partial_product_20(288) <= temp_mult_102(288);
partial_product_20(289) <= temp_mult_102(289);
partial_product_20(290) <= temp_mult_102(290);
partial_product_20(291) <= temp_mult_102(291);
partial_product_20(292) <= temp_mult_102(292);
partial_product_20(293) <= temp_mult_102(293);
partial_product_20(294) <= temp_mult_102(294);
partial_product_20(295) <= temp_mult_102(295);
partial_product_20(296) <= temp_mult_102(296);
partial_product_20(297) <= temp_mult_102(297);
partial_product_20(298) <= temp_mult_102(298);
partial_product_20(299) <= temp_mult_102(299);
partial_product_20(300) <= temp_mult_102(300);
partial_product_20(301) <= temp_mult_102(301);
partial_product_20(302) <= temp_mult_102(302);
partial_product_20(303) <= temp_mult_102(303);
partial_product_20(304) <= temp_mult_102(304);
partial_product_20(305) <= temp_mult_102(305);
partial_product_20(306) <= temp_mult_102(306);
partial_product_20(307) <= temp_mult_102(307);
partial_product_20(308) <= temp_mult_102(308);
partial_product_20(309) <= temp_mult_102(309);
partial_product_20(310) <= temp_mult_102(310);
partial_product_20(311) <= temp_mult_102(311);
partial_product_20(312) <= temp_mult_102(312);
partial_product_20(313) <= temp_mult_102(313);
partial_product_20(314) <= temp_mult_102(314);
partial_product_20(315) <= temp_mult_102(315);
partial_product_20(316) <= temp_mult_102(316);
partial_product_20(317) <= temp_mult_102(317);
partial_product_20(318) <= temp_mult_102(318);
partial_product_20(319) <= temp_mult_102(319);
partial_product_20(320) <= temp_mult_102(320);
partial_product_20(321) <= temp_mult_102(321);
partial_product_20(322) <= temp_mult_102(322);
partial_product_20(323) <= temp_mult_102(323);
partial_product_20(324) <= temp_mult_102(324);
partial_product_20(325) <= temp_mult_102(325);
partial_product_20(326) <= temp_mult_102(326);
partial_product_20(327) <= '0';
partial_product_20(328) <= '0';
partial_product_20(329) <= '0';
partial_product_20(330) <= '0';
partial_product_20(331) <= '0';
partial_product_20(332) <= '0';
partial_product_20(333) <= '0';
partial_product_20(334) <= '0';
partial_product_20(335) <= '0';
partial_product_20(336) <= '0';
partial_product_20(337) <= '0';
partial_product_20(338) <= '0';
partial_product_20(339) <= '0';
partial_product_20(340) <= '0';
partial_product_20(341) <= '0';
partial_product_20(342) <= '0';
partial_product_20(343) <= '0';
partial_product_20(344) <= '0';
partial_product_20(345) <= '0';
partial_product_20(346) <= '0';
partial_product_20(347) <= '0';
partial_product_20(348) <= '0';
partial_product_20(349) <= '0';
partial_product_20(350) <= '0';
partial_product_20(351) <= '0';
partial_product_20(352) <= '0';
partial_product_20(353) <= '0';
partial_product_20(354) <= '0';
partial_product_20(355) <= '0';
partial_product_20(356) <= '0';
partial_product_20(357) <= '0';
partial_product_20(358) <= '0';
partial_product_20(359) <= '0';
partial_product_20(360) <= '0';
partial_product_20(361) <= '0';
partial_product_20(362) <= '0';
partial_product_20(363) <= '0';
partial_product_20(364) <= '0';
partial_product_20(365) <= '0';
partial_product_20(366) <= '0';
partial_product_20(367) <= '0';
partial_product_20(368) <= '0';
partial_product_20(369) <= '0';
partial_product_20(370) <= '0';
partial_product_20(371) <= '0';
partial_product_20(372) <= '0';
partial_product_20(373) <= '0';
partial_product_20(374) <= '0';
partial_product_20(375) <= '0';
partial_product_20(376) <= '0';
partial_product_20(377) <= '0';
partial_product_20(378) <= '0';
partial_product_20(379) <= '0';
partial_product_20(380) <= '0';
partial_product_20(381) <= '0';
partial_product_20(382) <= '0';
partial_product_20(383) <= '0';
partial_product_20(384) <= '0';
partial_product_20(385) <= '0';
partial_product_20(386) <= '0';
partial_product_20(387) <= '0';
partial_product_20(388) <= '0';
partial_product_20(389) <= '0';
partial_product_20(390) <= '0';
partial_product_20(391) <= '0';
partial_product_20(392) <= '0';
partial_product_20(393) <= '0';
partial_product_20(394) <= '0';
partial_product_20(395) <= '0';
partial_product_20(396) <= '0';
partial_product_20(397) <= '0';
partial_product_20(398) <= '0';
partial_product_20(399) <= '0';
partial_product_20(400) <= '0';
partial_product_20(401) <= '0';
partial_product_20(402) <= '0';
partial_product_20(403) <= '0';
partial_product_20(404) <= '0';
partial_product_20(405) <= '0';
partial_product_20(406) <= '0';
partial_product_20(407) <= '0';
partial_product_20(408) <= '0';
partial_product_20(409) <= '0';
partial_product_20(410) <= '0';
partial_product_20(411) <= '0';
partial_product_20(412) <= '0';
partial_product_20(413) <= '0';
partial_product_20(414) <= '0';
partial_product_20(415) <= '0';
partial_product_20(416) <= '0';
partial_product_20(417) <= '0';
partial_product_20(418) <= '0';
partial_product_20(419) <= '0';
partial_product_20(420) <= '0';
partial_product_20(421) <= '0';
partial_product_20(422) <= '0';
partial_product_20(423) <= '0';
partial_product_20(424) <= '0';
partial_product_20(425) <= '0';
partial_product_20(426) <= '0';
partial_product_20(427) <= '0';
partial_product_20(428) <= '0';
partial_product_20(429) <= '0';
partial_product_20(430) <= '0';
partial_product_20(431) <= '0';
partial_product_20(432) <= '0';
partial_product_20(433) <= '0';
partial_product_20(434) <= '0';
partial_product_20(435) <= '0';
partial_product_20(436) <= '0';
partial_product_20(437) <= '0';
partial_product_20(438) <= '0';
partial_product_20(439) <= '0';
partial_product_20(440) <= '0';
partial_product_20(441) <= '0';
partial_product_20(442) <= '0';
partial_product_20(443) <= '0';
partial_product_20(444) <= '0';
partial_product_20(445) <= '0';
partial_product_20(446) <= '0';
partial_product_20(447) <= '0';
partial_product_20(448) <= '0';
partial_product_20(449) <= '0';
partial_product_20(450) <= '0';
partial_product_20(451) <= '0';
partial_product_20(452) <= '0';
partial_product_20(453) <= '0';
partial_product_20(454) <= '0';
partial_product_20(455) <= '0';
partial_product_20(456) <= '0';
partial_product_20(457) <= '0';
partial_product_20(458) <= '0';
partial_product_20(459) <= '0';
partial_product_20(460) <= '0';
partial_product_20(461) <= '0';
partial_product_20(462) <= '0';
partial_product_20(463) <= '0';
partial_product_20(464) <= '0';
partial_product_20(465) <= '0';
partial_product_20(466) <= '0';
partial_product_20(467) <= '0';
partial_product_20(468) <= '0';
partial_product_20(469) <= '0';
partial_product_20(470) <= '0';
partial_product_20(471) <= '0';
partial_product_20(472) <= '0';
partial_product_20(473) <= '0';
partial_product_20(474) <= '0';
partial_product_20(475) <= '0';
partial_product_20(476) <= '0';
partial_product_20(477) <= '0';
partial_product_20(478) <= '0';
partial_product_20(479) <= '0';
partial_product_20(480) <= '0';
partial_product_20(481) <= '0';
partial_product_20(482) <= '0';
partial_product_20(483) <= '0';
partial_product_20(484) <= '0';
partial_product_20(485) <= '0';
partial_product_20(486) <= '0';
partial_product_20(487) <= '0';
partial_product_20(488) <= '0';
partial_product_20(489) <= '0';
partial_product_20(490) <= '0';
partial_product_20(491) <= '0';
partial_product_20(492) <= '0';
partial_product_20(493) <= '0';
partial_product_20(494) <= '0';
partial_product_20(495) <= '0';
partial_product_20(496) <= '0';
partial_product_20(497) <= '0';
partial_product_20(498) <= '0';
partial_product_20(499) <= '0';
partial_product_20(500) <= '0';
partial_product_20(501) <= '0';
partial_product_20(502) <= '0';
partial_product_20(503) <= '0';
partial_product_20(504) <= '0';
partial_product_20(505) <= '0';
partial_product_20(506) <= '0';
partial_product_20(507) <= '0';
partial_product_20(508) <= '0';
partial_product_20(509) <= '0';
partial_product_20(510) <= '0';
partial_product_20(511) <= '0';
partial_product_20(512) <= '0';
partial_product_21(0) <= '0';
partial_product_21(1) <= '0';
partial_product_21(2) <= '0';
partial_product_21(3) <= '0';
partial_product_21(4) <= '0';
partial_product_21(5) <= '0';
partial_product_21(6) <= '0';
partial_product_21(7) <= '0';
partial_product_21(8) <= '0';
partial_product_21(9) <= '0';
partial_product_21(10) <= '0';
partial_product_21(11) <= '0';
partial_product_21(12) <= '0';
partial_product_21(13) <= '0';
partial_product_21(14) <= '0';
partial_product_21(15) <= '0';
partial_product_21(16) <= '0';
partial_product_21(17) <= '0';
partial_product_21(18) <= '0';
partial_product_21(19) <= '0';
partial_product_21(20) <= '0';
partial_product_21(21) <= '0';
partial_product_21(22) <= '0';
partial_product_21(23) <= '0';
partial_product_21(24) <= '0';
partial_product_21(25) <= '0';
partial_product_21(26) <= '0';
partial_product_21(27) <= '0';
partial_product_21(28) <= '0';
partial_product_21(29) <= '0';
partial_product_21(30) <= '0';
partial_product_21(31) <= '0';
partial_product_21(32) <= '0';
partial_product_21(33) <= '0';
partial_product_21(34) <= '0';
partial_product_21(35) <= '0';
partial_product_21(36) <= '0';
partial_product_21(37) <= '0';
partial_product_21(38) <= '0';
partial_product_21(39) <= '0';
partial_product_21(40) <= '0';
partial_product_21(41) <= '0';
partial_product_21(42) <= '0';
partial_product_21(43) <= '0';
partial_product_21(44) <= '0';
partial_product_21(45) <= '0';
partial_product_21(46) <= '0';
partial_product_21(47) <= '0';
partial_product_21(48) <= '0';
partial_product_21(49) <= '0';
partial_product_21(50) <= '0';
partial_product_21(51) <= '0';
partial_product_21(52) <= '0';
partial_product_21(53) <= '0';
partial_product_21(54) <= '0';
partial_product_21(55) <= '0';
partial_product_21(56) <= '0';
partial_product_21(57) <= '0';
partial_product_21(58) <= '0';
partial_product_21(59) <= '0';
partial_product_21(60) <= '0';
partial_product_21(61) <= '0';
partial_product_21(62) <= '0';
partial_product_21(63) <= '0';
partial_product_21(64) <= '0';
partial_product_21(65) <= '0';
partial_product_21(66) <= '0';
partial_product_21(67) <= '0';
partial_product_21(68) <= '0';
partial_product_21(69) <= '0';
partial_product_21(70) <= '0';
partial_product_21(71) <= '0';
partial_product_21(72) <= '0';
partial_product_21(73) <= '0';
partial_product_21(74) <= '0';
partial_product_21(75) <= '0';
partial_product_21(76) <= '0';
partial_product_21(77) <= '0';
partial_product_21(78) <= '0';
partial_product_21(79) <= '0';
partial_product_21(80) <= '0';
partial_product_21(81) <= '0';
partial_product_21(82) <= '0';
partial_product_21(83) <= '0';
partial_product_21(84) <= '0';
partial_product_21(85) <= '0';
partial_product_21(86) <= '0';
partial_product_21(87) <= '0';
partial_product_21(88) <= '0';
partial_product_21(89) <= '0';
partial_product_21(90) <= '0';
partial_product_21(91) <= '0';
partial_product_21(92) <= '0';
partial_product_21(93) <= '0';
partial_product_21(94) <= '0';
partial_product_21(95) <= '0';
partial_product_21(96) <= '0';
partial_product_21(97) <= '0';
partial_product_21(98) <= '0';
partial_product_21(99) <= '0';
partial_product_21(100) <= '0';
partial_product_21(101) <= '0';
partial_product_21(102) <= '0';
partial_product_21(103) <= '0';
partial_product_21(104) <= '0';
partial_product_21(105) <= '0';
partial_product_21(106) <= '0';
partial_product_21(107) <= '0';
partial_product_21(108) <= '0';
partial_product_21(109) <= '0';
partial_product_21(110) <= '0';
partial_product_21(111) <= '0';
partial_product_21(112) <= '0';
partial_product_21(113) <= '0';
partial_product_21(114) <= '0';
partial_product_21(115) <= '0';
partial_product_21(116) <= '0';
partial_product_21(117) <= '0';
partial_product_21(118) <= '0';
partial_product_21(119) <= '0';
partial_product_21(120) <= '0';
partial_product_21(121) <= '0';
partial_product_21(122) <= '0';
partial_product_21(123) <= '0';
partial_product_21(124) <= '0';
partial_product_21(125) <= '0';
partial_product_21(126) <= '0';
partial_product_21(127) <= '0';
partial_product_21(128) <= '0';
partial_product_21(129) <= '0';
partial_product_21(130) <= '0';
partial_product_21(131) <= '0';
partial_product_21(132) <= '0';
partial_product_21(133) <= '0';
partial_product_21(134) <= '0';
partial_product_21(135) <= '0';
partial_product_21(136) <= '0';
partial_product_21(137) <= '0';
partial_product_21(138) <= '0';
partial_product_21(139) <= '0';
partial_product_21(140) <= '0';
partial_product_21(141) <= '0';
partial_product_21(142) <= '0';
partial_product_21(143) <= '0';
partial_product_21(144) <= '0';
partial_product_21(145) <= '0';
partial_product_21(146) <= '0';
partial_product_21(147) <= '0';
partial_product_21(148) <= '0';
partial_product_21(149) <= '0';
partial_product_21(150) <= '0';
partial_product_21(151) <= '0';
partial_product_21(152) <= '0';
partial_product_21(153) <= '0';
partial_product_21(154) <= '0';
partial_product_21(155) <= '0';
partial_product_21(156) <= '0';
partial_product_21(157) <= '0';
partial_product_21(158) <= '0';
partial_product_21(159) <= '0';
partial_product_21(160) <= '0';
partial_product_21(161) <= '0';
partial_product_21(162) <= '0';
partial_product_21(163) <= '0';
partial_product_21(164) <= '0';
partial_product_21(165) <= '0';
partial_product_21(166) <= '0';
partial_product_21(167) <= '0';
partial_product_21(168) <= '0';
partial_product_21(169) <= '0';
partial_product_21(170) <= '0';
partial_product_21(171) <= '0';
partial_product_21(172) <= '0';
partial_product_21(173) <= '0';
partial_product_21(174) <= '0';
partial_product_21(175) <= '0';
partial_product_21(176) <= '0';
partial_product_21(177) <= '0';
partial_product_21(178) <= '0';
partial_product_21(179) <= '0';
partial_product_21(180) <= '0';
partial_product_21(181) <= '0';
partial_product_21(182) <= '0';
partial_product_21(183) <= '0';
partial_product_21(184) <= '0';
partial_product_21(185) <= '0';
partial_product_21(186) <= '0';
partial_product_21(187) <= '0';
partial_product_21(188) <= '0';
partial_product_21(189) <= '0';
partial_product_21(190) <= '0';
partial_product_21(191) <= '0';
partial_product_21(192) <= '0';
partial_product_21(193) <= '0';
partial_product_21(194) <= '0';
partial_product_21(195) <= '0';
partial_product_21(196) <= '0';
partial_product_21(197) <= '0';
partial_product_21(198) <= '0';
partial_product_21(199) <= '0';
partial_product_21(200) <= '0';
partial_product_21(201) <= '0';
partial_product_21(202) <= '0';
partial_product_21(203) <= '0';
partial_product_21(204) <= '0';
partial_product_21(205) <= '0';
partial_product_21(206) <= '0';
partial_product_21(207) <= '0';
partial_product_21(208) <= '0';
partial_product_21(209) <= '0';
partial_product_21(210) <= '0';
partial_product_21(211) <= '0';
partial_product_21(212) <= '0';
partial_product_21(213) <= '0';
partial_product_21(214) <= '0';
partial_product_21(215) <= '0';
partial_product_21(216) <= temp_mult_72(216);
partial_product_21(217) <= temp_mult_72(217);
partial_product_21(218) <= temp_mult_72(218);
partial_product_21(219) <= temp_mult_72(219);
partial_product_21(220) <= temp_mult_72(220);
partial_product_21(221) <= temp_mult_72(221);
partial_product_21(222) <= temp_mult_72(222);
partial_product_21(223) <= temp_mult_72(223);
partial_product_21(224) <= temp_mult_72(224);
partial_product_21(225) <= temp_mult_72(225);
partial_product_21(226) <= temp_mult_72(226);
partial_product_21(227) <= temp_mult_72(227);
partial_product_21(228) <= temp_mult_72(228);
partial_product_21(229) <= temp_mult_72(229);
partial_product_21(230) <= temp_mult_72(230);
partial_product_21(231) <= temp_mult_72(231);
partial_product_21(232) <= temp_mult_72(232);
partial_product_21(233) <= temp_mult_72(233);
partial_product_21(234) <= temp_mult_72(234);
partial_product_21(235) <= temp_mult_72(235);
partial_product_21(236) <= temp_mult_72(236);
partial_product_21(237) <= temp_mult_72(237);
partial_product_21(238) <= temp_mult_72(238);
partial_product_21(239) <= temp_mult_72(239);
partial_product_21(240) <= temp_mult_72(240);
partial_product_21(241) <= temp_mult_72(241);
partial_product_21(242) <= temp_mult_72(242);
partial_product_21(243) <= temp_mult_72(243);
partial_product_21(244) <= temp_mult_72(244);
partial_product_21(245) <= temp_mult_72(245);
partial_product_21(246) <= temp_mult_72(246);
partial_product_21(247) <= temp_mult_72(247);
partial_product_21(248) <= temp_mult_72(248);
partial_product_21(249) <= temp_mult_72(249);
partial_product_21(250) <= temp_mult_72(250);
partial_product_21(251) <= temp_mult_72(251);
partial_product_21(252) <= temp_mult_72(252);
partial_product_21(253) <= temp_mult_72(253);
partial_product_21(254) <= temp_mult_72(254);
partial_product_21(255) <= temp_mult_72(255);
partial_product_21(256) <= temp_mult_72(256);
partial_product_21(257) <= '0';
partial_product_21(258) <= '0';
partial_product_21(259) <= '0';
partial_product_21(260) <= '0';
partial_product_21(261) <= '0';
partial_product_21(262) <= temp_mult_94(262);
partial_product_21(263) <= temp_mult_94(263);
partial_product_21(264) <= temp_mult_94(264);
partial_product_21(265) <= temp_mult_94(265);
partial_product_21(266) <= temp_mult_94(266);
partial_product_21(267) <= temp_mult_94(267);
partial_product_21(268) <= temp_mult_94(268);
partial_product_21(269) <= temp_mult_94(269);
partial_product_21(270) <= temp_mult_94(270);
partial_product_21(271) <= temp_mult_94(271);
partial_product_21(272) <= temp_mult_94(272);
partial_product_21(273) <= temp_mult_94(273);
partial_product_21(274) <= temp_mult_94(274);
partial_product_21(275) <= temp_mult_94(275);
partial_product_21(276) <= temp_mult_94(276);
partial_product_21(277) <= temp_mult_94(277);
partial_product_21(278) <= temp_mult_94(278);
partial_product_21(279) <= temp_mult_94(279);
partial_product_21(280) <= temp_mult_94(280);
partial_product_21(281) <= temp_mult_94(281);
partial_product_21(282) <= temp_mult_94(282);
partial_product_21(283) <= temp_mult_94(283);
partial_product_21(284) <= temp_mult_94(284);
partial_product_21(285) <= temp_mult_94(285);
partial_product_21(286) <= temp_mult_94(286);
partial_product_21(287) <= temp_mult_94(287);
partial_product_21(288) <= temp_mult_94(288);
partial_product_21(289) <= temp_mult_94(289);
partial_product_21(290) <= temp_mult_94(290);
partial_product_21(291) <= temp_mult_94(291);
partial_product_21(292) <= temp_mult_94(292);
partial_product_21(293) <= temp_mult_94(293);
partial_product_21(294) <= temp_mult_94(294);
partial_product_21(295) <= temp_mult_94(295);
partial_product_21(296) <= temp_mult_94(296);
partial_product_21(297) <= temp_mult_94(297);
partial_product_21(298) <= temp_mult_94(298);
partial_product_21(299) <= temp_mult_94(299);
partial_product_21(300) <= temp_mult_94(300);
partial_product_21(301) <= temp_mult_94(301);
partial_product_21(302) <= temp_mult_94(302);
partial_product_21(303) <= '0';
partial_product_21(304) <= '0';
partial_product_21(305) <= '0';
partial_product_21(306) <= '0';
partial_product_21(307) <= '0';
partial_product_21(308) <= '0';
partial_product_21(309) <= '0';
partial_product_21(310) <= '0';
partial_product_21(311) <= '0';
partial_product_21(312) <= '0';
partial_product_21(313) <= '0';
partial_product_21(314) <= '0';
partial_product_21(315) <= '0';
partial_product_21(316) <= '0';
partial_product_21(317) <= '0';
partial_product_21(318) <= '0';
partial_product_21(319) <= '0';
partial_product_21(320) <= '0';
partial_product_21(321) <= '0';
partial_product_21(322) <= '0';
partial_product_21(323) <= '0';
partial_product_21(324) <= '0';
partial_product_21(325) <= '0';
partial_product_21(326) <= '0';
partial_product_21(327) <= '0';
partial_product_21(328) <= '0';
partial_product_21(329) <= '0';
partial_product_21(330) <= '0';
partial_product_21(331) <= '0';
partial_product_21(332) <= '0';
partial_product_21(333) <= '0';
partial_product_21(334) <= '0';
partial_product_21(335) <= '0';
partial_product_21(336) <= '0';
partial_product_21(337) <= '0';
partial_product_21(338) <= '0';
partial_product_21(339) <= '0';
partial_product_21(340) <= '0';
partial_product_21(341) <= '0';
partial_product_21(342) <= '0';
partial_product_21(343) <= '0';
partial_product_21(344) <= '0';
partial_product_21(345) <= '0';
partial_product_21(346) <= '0';
partial_product_21(347) <= '0';
partial_product_21(348) <= '0';
partial_product_21(349) <= '0';
partial_product_21(350) <= '0';
partial_product_21(351) <= '0';
partial_product_21(352) <= '0';
partial_product_21(353) <= '0';
partial_product_21(354) <= '0';
partial_product_21(355) <= '0';
partial_product_21(356) <= '0';
partial_product_21(357) <= '0';
partial_product_21(358) <= '0';
partial_product_21(359) <= '0';
partial_product_21(360) <= '0';
partial_product_21(361) <= '0';
partial_product_21(362) <= '0';
partial_product_21(363) <= '0';
partial_product_21(364) <= '0';
partial_product_21(365) <= '0';
partial_product_21(366) <= '0';
partial_product_21(367) <= '0';
partial_product_21(368) <= '0';
partial_product_21(369) <= '0';
partial_product_21(370) <= '0';
partial_product_21(371) <= '0';
partial_product_21(372) <= '0';
partial_product_21(373) <= '0';
partial_product_21(374) <= '0';
partial_product_21(375) <= '0';
partial_product_21(376) <= '0';
partial_product_21(377) <= '0';
partial_product_21(378) <= '0';
partial_product_21(379) <= '0';
partial_product_21(380) <= '0';
partial_product_21(381) <= '0';
partial_product_21(382) <= '0';
partial_product_21(383) <= '0';
partial_product_21(384) <= '0';
partial_product_21(385) <= '0';
partial_product_21(386) <= '0';
partial_product_21(387) <= '0';
partial_product_21(388) <= '0';
partial_product_21(389) <= '0';
partial_product_21(390) <= '0';
partial_product_21(391) <= '0';
partial_product_21(392) <= '0';
partial_product_21(393) <= '0';
partial_product_21(394) <= '0';
partial_product_21(395) <= '0';
partial_product_21(396) <= '0';
partial_product_21(397) <= '0';
partial_product_21(398) <= '0';
partial_product_21(399) <= '0';
partial_product_21(400) <= '0';
partial_product_21(401) <= '0';
partial_product_21(402) <= '0';
partial_product_21(403) <= '0';
partial_product_21(404) <= '0';
partial_product_21(405) <= '0';
partial_product_21(406) <= '0';
partial_product_21(407) <= '0';
partial_product_21(408) <= '0';
partial_product_21(409) <= '0';
partial_product_21(410) <= '0';
partial_product_21(411) <= '0';
partial_product_21(412) <= '0';
partial_product_21(413) <= '0';
partial_product_21(414) <= '0';
partial_product_21(415) <= '0';
partial_product_21(416) <= '0';
partial_product_21(417) <= '0';
partial_product_21(418) <= '0';
partial_product_21(419) <= '0';
partial_product_21(420) <= '0';
partial_product_21(421) <= '0';
partial_product_21(422) <= '0';
partial_product_21(423) <= '0';
partial_product_21(424) <= '0';
partial_product_21(425) <= '0';
partial_product_21(426) <= '0';
partial_product_21(427) <= '0';
partial_product_21(428) <= '0';
partial_product_21(429) <= '0';
partial_product_21(430) <= '0';
partial_product_21(431) <= '0';
partial_product_21(432) <= '0';
partial_product_21(433) <= '0';
partial_product_21(434) <= '0';
partial_product_21(435) <= '0';
partial_product_21(436) <= '0';
partial_product_21(437) <= '0';
partial_product_21(438) <= '0';
partial_product_21(439) <= '0';
partial_product_21(440) <= '0';
partial_product_21(441) <= '0';
partial_product_21(442) <= '0';
partial_product_21(443) <= '0';
partial_product_21(444) <= '0';
partial_product_21(445) <= '0';
partial_product_21(446) <= '0';
partial_product_21(447) <= '0';
partial_product_21(448) <= '0';
partial_product_21(449) <= '0';
partial_product_21(450) <= '0';
partial_product_21(451) <= '0';
partial_product_21(452) <= '0';
partial_product_21(453) <= '0';
partial_product_21(454) <= '0';
partial_product_21(455) <= '0';
partial_product_21(456) <= '0';
partial_product_21(457) <= '0';
partial_product_21(458) <= '0';
partial_product_21(459) <= '0';
partial_product_21(460) <= '0';
partial_product_21(461) <= '0';
partial_product_21(462) <= '0';
partial_product_21(463) <= '0';
partial_product_21(464) <= '0';
partial_product_21(465) <= '0';
partial_product_21(466) <= '0';
partial_product_21(467) <= '0';
partial_product_21(468) <= '0';
partial_product_21(469) <= '0';
partial_product_21(470) <= '0';
partial_product_21(471) <= '0';
partial_product_21(472) <= '0';
partial_product_21(473) <= '0';
partial_product_21(474) <= '0';
partial_product_21(475) <= '0';
partial_product_21(476) <= '0';
partial_product_21(477) <= '0';
partial_product_21(478) <= '0';
partial_product_21(479) <= '0';
partial_product_21(480) <= '0';
partial_product_21(481) <= '0';
partial_product_21(482) <= '0';
partial_product_21(483) <= '0';
partial_product_21(484) <= '0';
partial_product_21(485) <= '0';
partial_product_21(486) <= '0';
partial_product_21(487) <= '0';
partial_product_21(488) <= '0';
partial_product_21(489) <= '0';
partial_product_21(490) <= '0';
partial_product_21(491) <= '0';
partial_product_21(492) <= '0';
partial_product_21(493) <= '0';
partial_product_21(494) <= '0';
partial_product_21(495) <= '0';
partial_product_21(496) <= '0';
partial_product_21(497) <= '0';
partial_product_21(498) <= '0';
partial_product_21(499) <= '0';
partial_product_21(500) <= '0';
partial_product_21(501) <= '0';
partial_product_21(502) <= '0';
partial_product_21(503) <= '0';
partial_product_21(504) <= '0';
partial_product_21(505) <= '0';
partial_product_21(506) <= '0';
partial_product_21(507) <= '0';
partial_product_21(508) <= '0';
partial_product_21(509) <= '0';
partial_product_21(510) <= '0';
partial_product_21(511) <= '0';
partial_product_21(512) <= '0';
partial_product_22(0) <= '0';
partial_product_22(1) <= '0';
partial_product_22(2) <= '0';
partial_product_22(3) <= '0';
partial_product_22(4) <= '0';
partial_product_22(5) <= '0';
partial_product_22(6) <= '0';
partial_product_22(7) <= '0';
partial_product_22(8) <= '0';
partial_product_22(9) <= '0';
partial_product_22(10) <= '0';
partial_product_22(11) <= '0';
partial_product_22(12) <= '0';
partial_product_22(13) <= '0';
partial_product_22(14) <= '0';
partial_product_22(15) <= '0';
partial_product_22(16) <= '0';
partial_product_22(17) <= '0';
partial_product_22(18) <= '0';
partial_product_22(19) <= '0';
partial_product_22(20) <= '0';
partial_product_22(21) <= '0';
partial_product_22(22) <= '0';
partial_product_22(23) <= '0';
partial_product_22(24) <= '0';
partial_product_22(25) <= '0';
partial_product_22(26) <= '0';
partial_product_22(27) <= '0';
partial_product_22(28) <= '0';
partial_product_22(29) <= '0';
partial_product_22(30) <= '0';
partial_product_22(31) <= '0';
partial_product_22(32) <= '0';
partial_product_22(33) <= '0';
partial_product_22(34) <= '0';
partial_product_22(35) <= '0';
partial_product_22(36) <= '0';
partial_product_22(37) <= '0';
partial_product_22(38) <= '0';
partial_product_22(39) <= '0';
partial_product_22(40) <= '0';
partial_product_22(41) <= '0';
partial_product_22(42) <= '0';
partial_product_22(43) <= '0';
partial_product_22(44) <= '0';
partial_product_22(45) <= '0';
partial_product_22(46) <= '0';
partial_product_22(47) <= '0';
partial_product_22(48) <= '0';
partial_product_22(49) <= '0';
partial_product_22(50) <= '0';
partial_product_22(51) <= '0';
partial_product_22(52) <= '0';
partial_product_22(53) <= '0';
partial_product_22(54) <= '0';
partial_product_22(55) <= '0';
partial_product_22(56) <= '0';
partial_product_22(57) <= '0';
partial_product_22(58) <= '0';
partial_product_22(59) <= '0';
partial_product_22(60) <= '0';
partial_product_22(61) <= '0';
partial_product_22(62) <= '0';
partial_product_22(63) <= '0';
partial_product_22(64) <= '0';
partial_product_22(65) <= '0';
partial_product_22(66) <= '0';
partial_product_22(67) <= '0';
partial_product_22(68) <= '0';
partial_product_22(69) <= '0';
partial_product_22(70) <= '0';
partial_product_22(71) <= '0';
partial_product_22(72) <= '0';
partial_product_22(73) <= '0';
partial_product_22(74) <= '0';
partial_product_22(75) <= '0';
partial_product_22(76) <= '0';
partial_product_22(77) <= '0';
partial_product_22(78) <= '0';
partial_product_22(79) <= '0';
partial_product_22(80) <= '0';
partial_product_22(81) <= '0';
partial_product_22(82) <= '0';
partial_product_22(83) <= '0';
partial_product_22(84) <= '0';
partial_product_22(85) <= '0';
partial_product_22(86) <= '0';
partial_product_22(87) <= '0';
partial_product_22(88) <= '0';
partial_product_22(89) <= '0';
partial_product_22(90) <= '0';
partial_product_22(91) <= '0';
partial_product_22(92) <= '0';
partial_product_22(93) <= '0';
partial_product_22(94) <= '0';
partial_product_22(95) <= '0';
partial_product_22(96) <= '0';
partial_product_22(97) <= '0';
partial_product_22(98) <= '0';
partial_product_22(99) <= '0';
partial_product_22(100) <= '0';
partial_product_22(101) <= '0';
partial_product_22(102) <= '0';
partial_product_22(103) <= '0';
partial_product_22(104) <= '0';
partial_product_22(105) <= '0';
partial_product_22(106) <= '0';
partial_product_22(107) <= '0';
partial_product_22(108) <= '0';
partial_product_22(109) <= '0';
partial_product_22(110) <= '0';
partial_product_22(111) <= '0';
partial_product_22(112) <= '0';
partial_product_22(113) <= '0';
partial_product_22(114) <= '0';
partial_product_22(115) <= '0';
partial_product_22(116) <= '0';
partial_product_22(117) <= '0';
partial_product_22(118) <= '0';
partial_product_22(119) <= '0';
partial_product_22(120) <= '0';
partial_product_22(121) <= '0';
partial_product_22(122) <= '0';
partial_product_22(123) <= '0';
partial_product_22(124) <= '0';
partial_product_22(125) <= '0';
partial_product_22(126) <= '0';
partial_product_22(127) <= '0';
partial_product_22(128) <= '0';
partial_product_22(129) <= '0';
partial_product_22(130) <= '0';
partial_product_22(131) <= '0';
partial_product_22(132) <= '0';
partial_product_22(133) <= '0';
partial_product_22(134) <= '0';
partial_product_22(135) <= '0';
partial_product_22(136) <= '0';
partial_product_22(137) <= '0';
partial_product_22(138) <= '0';
partial_product_22(139) <= '0';
partial_product_22(140) <= '0';
partial_product_22(141) <= '0';
partial_product_22(142) <= '0';
partial_product_22(143) <= '0';
partial_product_22(144) <= '0';
partial_product_22(145) <= '0';
partial_product_22(146) <= '0';
partial_product_22(147) <= '0';
partial_product_22(148) <= '0';
partial_product_22(149) <= '0';
partial_product_22(150) <= '0';
partial_product_22(151) <= '0';
partial_product_22(152) <= '0';
partial_product_22(153) <= '0';
partial_product_22(154) <= '0';
partial_product_22(155) <= '0';
partial_product_22(156) <= '0';
partial_product_22(157) <= '0';
partial_product_22(158) <= '0';
partial_product_22(159) <= '0';
partial_product_22(160) <= '0';
partial_product_22(161) <= '0';
partial_product_22(162) <= '0';
partial_product_22(163) <= '0';
partial_product_22(164) <= '0';
partial_product_22(165) <= '0';
partial_product_22(166) <= '0';
partial_product_22(167) <= '0';
partial_product_22(168) <= '0';
partial_product_22(169) <= '0';
partial_product_22(170) <= '0';
partial_product_22(171) <= '0';
partial_product_22(172) <= '0';
partial_product_22(173) <= '0';
partial_product_22(174) <= '0';
partial_product_22(175) <= '0';
partial_product_22(176) <= '0';
partial_product_22(177) <= '0';
partial_product_22(178) <= '0';
partial_product_22(179) <= '0';
partial_product_22(180) <= '0';
partial_product_22(181) <= '0';
partial_product_22(182) <= '0';
partial_product_22(183) <= '0';
partial_product_22(184) <= '0';
partial_product_22(185) <= '0';
partial_product_22(186) <= '0';
partial_product_22(187) <= '0';
partial_product_22(188) <= '0';
partial_product_22(189) <= '0';
partial_product_22(190) <= '0';
partial_product_22(191) <= '0';
partial_product_22(192) <= '0';
partial_product_22(193) <= '0';
partial_product_22(194) <= '0';
partial_product_22(195) <= '0';
partial_product_22(196) <= '0';
partial_product_22(197) <= '0';
partial_product_22(198) <= '0';
partial_product_22(199) <= '0';
partial_product_22(200) <= '0';
partial_product_22(201) <= '0';
partial_product_22(202) <= '0';
partial_product_22(203) <= '0';
partial_product_22(204) <= '0';
partial_product_22(205) <= '0';
partial_product_22(206) <= '0';
partial_product_22(207) <= '0';
partial_product_22(208) <= '0';
partial_product_22(209) <= '0';
partial_product_22(210) <= '0';
partial_product_22(211) <= '0';
partial_product_22(212) <= '0';
partial_product_22(213) <= '0';
partial_product_22(214) <= '0';
partial_product_22(215) <= '0';
partial_product_22(216) <= '0';
partial_product_22(217) <= '0';
partial_product_22(218) <= '0';
partial_product_22(219) <= '0';
partial_product_22(220) <= '0';
partial_product_22(221) <= temp_mult_85(221);
partial_product_22(222) <= temp_mult_85(222);
partial_product_22(223) <= temp_mult_85(223);
partial_product_22(224) <= temp_mult_85(224);
partial_product_22(225) <= temp_mult_85(225);
partial_product_22(226) <= temp_mult_85(226);
partial_product_22(227) <= temp_mult_85(227);
partial_product_22(228) <= temp_mult_85(228);
partial_product_22(229) <= temp_mult_85(229);
partial_product_22(230) <= temp_mult_85(230);
partial_product_22(231) <= temp_mult_85(231);
partial_product_22(232) <= temp_mult_85(232);
partial_product_22(233) <= temp_mult_85(233);
partial_product_22(234) <= temp_mult_85(234);
partial_product_22(235) <= temp_mult_85(235);
partial_product_22(236) <= temp_mult_85(236);
partial_product_22(237) <= temp_mult_85(237);
partial_product_22(238) <= temp_mult_85(238);
partial_product_22(239) <= temp_mult_85(239);
partial_product_22(240) <= temp_mult_85(240);
partial_product_22(241) <= temp_mult_85(241);
partial_product_22(242) <= temp_mult_85(242);
partial_product_22(243) <= temp_mult_85(243);
partial_product_22(244) <= temp_mult_85(244);
partial_product_22(245) <= temp_mult_85(245);
partial_product_22(246) <= temp_mult_85(246);
partial_product_22(247) <= temp_mult_85(247);
partial_product_22(248) <= temp_mult_85(248);
partial_product_22(249) <= temp_mult_85(249);
partial_product_22(250) <= temp_mult_85(250);
partial_product_22(251) <= temp_mult_85(251);
partial_product_22(252) <= temp_mult_85(252);
partial_product_22(253) <= temp_mult_85(253);
partial_product_22(254) <= temp_mult_85(254);
partial_product_22(255) <= temp_mult_85(255);
partial_product_22(256) <= temp_mult_85(256);
partial_product_22(257) <= temp_mult_85(257);
partial_product_22(258) <= temp_mult_85(258);
partial_product_22(259) <= temp_mult_85(259);
partial_product_22(260) <= temp_mult_85(260);
partial_product_22(261) <= temp_mult_85(261);
partial_product_22(262) <= '0';
partial_product_22(263) <= '0';
partial_product_22(264) <= '0';
partial_product_22(265) <= '0';
partial_product_22(266) <= '0';
partial_product_22(267) <= '0';
partial_product_22(268) <= '0';
partial_product_22(269) <= '0';
partial_product_22(270) <= '0';
partial_product_22(271) <= '0';
partial_product_22(272) <= '0';
partial_product_22(273) <= '0';
partial_product_22(274) <= '0';
partial_product_22(275) <= '0';
partial_product_22(276) <= '0';
partial_product_22(277) <= '0';
partial_product_22(278) <= '0';
partial_product_22(279) <= '0';
partial_product_22(280) <= '0';
partial_product_22(281) <= '0';
partial_product_22(282) <= '0';
partial_product_22(283) <= '0';
partial_product_22(284) <= '0';
partial_product_22(285) <= '0';
partial_product_22(286) <= '0';
partial_product_22(287) <= '0';
partial_product_22(288) <= '0';
partial_product_22(289) <= '0';
partial_product_22(290) <= '0';
partial_product_22(291) <= '0';
partial_product_22(292) <= '0';
partial_product_22(293) <= '0';
partial_product_22(294) <= '0';
partial_product_22(295) <= '0';
partial_product_22(296) <= '0';
partial_product_22(297) <= '0';
partial_product_22(298) <= '0';
partial_product_22(299) <= '0';
partial_product_22(300) <= '0';
partial_product_22(301) <= '0';
partial_product_22(302) <= '0';
partial_product_22(303) <= '0';
partial_product_22(304) <= '0';
partial_product_22(305) <= '0';
partial_product_22(306) <= '0';
partial_product_22(307) <= '0';
partial_product_22(308) <= '0';
partial_product_22(309) <= '0';
partial_product_22(310) <= '0';
partial_product_22(311) <= '0';
partial_product_22(312) <= '0';
partial_product_22(313) <= '0';
partial_product_22(314) <= '0';
partial_product_22(315) <= '0';
partial_product_22(316) <= '0';
partial_product_22(317) <= '0';
partial_product_22(318) <= '0';
partial_product_22(319) <= '0';
partial_product_22(320) <= '0';
partial_product_22(321) <= '0';
partial_product_22(322) <= '0';
partial_product_22(323) <= '0';
partial_product_22(324) <= '0';
partial_product_22(325) <= '0';
partial_product_22(326) <= '0';
partial_product_22(327) <= '0';
partial_product_22(328) <= '0';
partial_product_22(329) <= '0';
partial_product_22(330) <= '0';
partial_product_22(331) <= '0';
partial_product_22(332) <= '0';
partial_product_22(333) <= '0';
partial_product_22(334) <= '0';
partial_product_22(335) <= '0';
partial_product_22(336) <= '0';
partial_product_22(337) <= '0';
partial_product_22(338) <= '0';
partial_product_22(339) <= '0';
partial_product_22(340) <= '0';
partial_product_22(341) <= '0';
partial_product_22(342) <= '0';
partial_product_22(343) <= '0';
partial_product_22(344) <= '0';
partial_product_22(345) <= '0';
partial_product_22(346) <= '0';
partial_product_22(347) <= '0';
partial_product_22(348) <= '0';
partial_product_22(349) <= '0';
partial_product_22(350) <= '0';
partial_product_22(351) <= '0';
partial_product_22(352) <= '0';
partial_product_22(353) <= '0';
partial_product_22(354) <= '0';
partial_product_22(355) <= '0';
partial_product_22(356) <= '0';
partial_product_22(357) <= '0';
partial_product_22(358) <= '0';
partial_product_22(359) <= '0';
partial_product_22(360) <= '0';
partial_product_22(361) <= '0';
partial_product_22(362) <= '0';
partial_product_22(363) <= '0';
partial_product_22(364) <= '0';
partial_product_22(365) <= '0';
partial_product_22(366) <= '0';
partial_product_22(367) <= '0';
partial_product_22(368) <= '0';
partial_product_22(369) <= '0';
partial_product_22(370) <= '0';
partial_product_22(371) <= '0';
partial_product_22(372) <= '0';
partial_product_22(373) <= '0';
partial_product_22(374) <= '0';
partial_product_22(375) <= '0';
partial_product_22(376) <= '0';
partial_product_22(377) <= '0';
partial_product_22(378) <= '0';
partial_product_22(379) <= '0';
partial_product_22(380) <= '0';
partial_product_22(381) <= '0';
partial_product_22(382) <= '0';
partial_product_22(383) <= '0';
partial_product_22(384) <= '0';
partial_product_22(385) <= '0';
partial_product_22(386) <= '0';
partial_product_22(387) <= '0';
partial_product_22(388) <= '0';
partial_product_22(389) <= '0';
partial_product_22(390) <= '0';
partial_product_22(391) <= '0';
partial_product_22(392) <= '0';
partial_product_22(393) <= '0';
partial_product_22(394) <= '0';
partial_product_22(395) <= '0';
partial_product_22(396) <= '0';
partial_product_22(397) <= '0';
partial_product_22(398) <= '0';
partial_product_22(399) <= '0';
partial_product_22(400) <= '0';
partial_product_22(401) <= '0';
partial_product_22(402) <= '0';
partial_product_22(403) <= '0';
partial_product_22(404) <= '0';
partial_product_22(405) <= '0';
partial_product_22(406) <= '0';
partial_product_22(407) <= '0';
partial_product_22(408) <= '0';
partial_product_22(409) <= '0';
partial_product_22(410) <= '0';
partial_product_22(411) <= '0';
partial_product_22(412) <= '0';
partial_product_22(413) <= '0';
partial_product_22(414) <= '0';
partial_product_22(415) <= '0';
partial_product_22(416) <= '0';
partial_product_22(417) <= '0';
partial_product_22(418) <= '0';
partial_product_22(419) <= '0';
partial_product_22(420) <= '0';
partial_product_22(421) <= '0';
partial_product_22(422) <= '0';
partial_product_22(423) <= '0';
partial_product_22(424) <= '0';
partial_product_22(425) <= '0';
partial_product_22(426) <= '0';
partial_product_22(427) <= '0';
partial_product_22(428) <= '0';
partial_product_22(429) <= '0';
partial_product_22(430) <= '0';
partial_product_22(431) <= '0';
partial_product_22(432) <= '0';
partial_product_22(433) <= '0';
partial_product_22(434) <= '0';
partial_product_22(435) <= '0';
partial_product_22(436) <= '0';
partial_product_22(437) <= '0';
partial_product_22(438) <= '0';
partial_product_22(439) <= '0';
partial_product_22(440) <= '0';
partial_product_22(441) <= '0';
partial_product_22(442) <= '0';
partial_product_22(443) <= '0';
partial_product_22(444) <= '0';
partial_product_22(445) <= '0';
partial_product_22(446) <= '0';
partial_product_22(447) <= '0';
partial_product_22(448) <= '0';
partial_product_22(449) <= '0';
partial_product_22(450) <= '0';
partial_product_22(451) <= '0';
partial_product_22(452) <= '0';
partial_product_22(453) <= '0';
partial_product_22(454) <= '0';
partial_product_22(455) <= '0';
partial_product_22(456) <= '0';
partial_product_22(457) <= '0';
partial_product_22(458) <= '0';
partial_product_22(459) <= '0';
partial_product_22(460) <= '0';
partial_product_22(461) <= '0';
partial_product_22(462) <= '0';
partial_product_22(463) <= '0';
partial_product_22(464) <= '0';
partial_product_22(465) <= '0';
partial_product_22(466) <= '0';
partial_product_22(467) <= '0';
partial_product_22(468) <= '0';
partial_product_22(469) <= '0';
partial_product_22(470) <= '0';
partial_product_22(471) <= '0';
partial_product_22(472) <= '0';
partial_product_22(473) <= '0';
partial_product_22(474) <= '0';
partial_product_22(475) <= '0';
partial_product_22(476) <= '0';
partial_product_22(477) <= '0';
partial_product_22(478) <= '0';
partial_product_22(479) <= '0';
partial_product_22(480) <= '0';
partial_product_22(481) <= '0';
partial_product_22(482) <= '0';
partial_product_22(483) <= '0';
partial_product_22(484) <= '0';
partial_product_22(485) <= '0';
partial_product_22(486) <= '0';
partial_product_22(487) <= '0';
partial_product_22(488) <= '0';
partial_product_22(489) <= '0';
partial_product_22(490) <= '0';
partial_product_22(491) <= '0';
partial_product_22(492) <= '0';
partial_product_22(493) <= '0';
partial_product_22(494) <= '0';
partial_product_22(495) <= '0';
partial_product_22(496) <= '0';
partial_product_22(497) <= '0';
partial_product_22(498) <= '0';
partial_product_22(499) <= '0';
partial_product_22(500) <= '0';
partial_product_22(501) <= '0';
partial_product_22(502) <= '0';
partial_product_22(503) <= '0';
partial_product_22(504) <= '0';
partial_product_22(505) <= '0';
partial_product_22(506) <= '0';
partial_product_22(507) <= '0';
partial_product_22(508) <= '0';
partial_product_22(509) <= '0';
partial_product_22(510) <= '0';
partial_product_22(511) <= '0';
partial_product_22(512) <= '0';
partial_product_23(0) <= '0';
partial_product_23(1) <= '0';
partial_product_23(2) <= '0';
partial_product_23(3) <= '0';
partial_product_23(4) <= '0';
partial_product_23(5) <= '0';
partial_product_23(6) <= '0';
partial_product_23(7) <= '0';
partial_product_23(8) <= '0';
partial_product_23(9) <= '0';
partial_product_23(10) <= '0';
partial_product_23(11) <= '0';
partial_product_23(12) <= '0';
partial_product_23(13) <= '0';
partial_product_23(14) <= '0';
partial_product_23(15) <= '0';
partial_product_23(16) <= '0';
partial_product_23(17) <= '0';
partial_product_23(18) <= '0';
partial_product_23(19) <= '0';
partial_product_23(20) <= '0';
partial_product_23(21) <= '0';
partial_product_23(22) <= '0';
partial_product_23(23) <= '0';
partial_product_23(24) <= '0';
partial_product_23(25) <= '0';
partial_product_23(26) <= '0';
partial_product_23(27) <= '0';
partial_product_23(28) <= '0';
partial_product_23(29) <= '0';
partial_product_23(30) <= '0';
partial_product_23(31) <= '0';
partial_product_23(32) <= '0';
partial_product_23(33) <= '0';
partial_product_23(34) <= '0';
partial_product_23(35) <= '0';
partial_product_23(36) <= '0';
partial_product_23(37) <= '0';
partial_product_23(38) <= '0';
partial_product_23(39) <= '0';
partial_product_23(40) <= '0';
partial_product_23(41) <= '0';
partial_product_23(42) <= '0';
partial_product_23(43) <= '0';
partial_product_23(44) <= '0';
partial_product_23(45) <= '0';
partial_product_23(46) <= '0';
partial_product_23(47) <= '0';
partial_product_23(48) <= '0';
partial_product_23(49) <= '0';
partial_product_23(50) <= '0';
partial_product_23(51) <= '0';
partial_product_23(52) <= '0';
partial_product_23(53) <= '0';
partial_product_23(54) <= '0';
partial_product_23(55) <= '0';
partial_product_23(56) <= '0';
partial_product_23(57) <= '0';
partial_product_23(58) <= '0';
partial_product_23(59) <= '0';
partial_product_23(60) <= '0';
partial_product_23(61) <= '0';
partial_product_23(62) <= '0';
partial_product_23(63) <= '0';
partial_product_23(64) <= '0';
partial_product_23(65) <= '0';
partial_product_23(66) <= '0';
partial_product_23(67) <= '0';
partial_product_23(68) <= '0';
partial_product_23(69) <= '0';
partial_product_23(70) <= '0';
partial_product_23(71) <= '0';
partial_product_23(72) <= '0';
partial_product_23(73) <= '0';
partial_product_23(74) <= '0';
partial_product_23(75) <= '0';
partial_product_23(76) <= '0';
partial_product_23(77) <= '0';
partial_product_23(78) <= '0';
partial_product_23(79) <= '0';
partial_product_23(80) <= '0';
partial_product_23(81) <= '0';
partial_product_23(82) <= '0';
partial_product_23(83) <= '0';
partial_product_23(84) <= '0';
partial_product_23(85) <= '0';
partial_product_23(86) <= '0';
partial_product_23(87) <= '0';
partial_product_23(88) <= '0';
partial_product_23(89) <= '0';
partial_product_23(90) <= '0';
partial_product_23(91) <= '0';
partial_product_23(92) <= '0';
partial_product_23(93) <= '0';
partial_product_23(94) <= '0';
partial_product_23(95) <= '0';
partial_product_23(96) <= '0';
partial_product_23(97) <= '0';
partial_product_23(98) <= '0';
partial_product_23(99) <= '0';
partial_product_23(100) <= '0';
partial_product_23(101) <= '0';
partial_product_23(102) <= '0';
partial_product_23(103) <= '0';
partial_product_23(104) <= '0';
partial_product_23(105) <= '0';
partial_product_23(106) <= '0';
partial_product_23(107) <= '0';
partial_product_23(108) <= '0';
partial_product_23(109) <= '0';
partial_product_23(110) <= '0';
partial_product_23(111) <= '0';
partial_product_23(112) <= '0';
partial_product_23(113) <= '0';
partial_product_23(114) <= '0';
partial_product_23(115) <= '0';
partial_product_23(116) <= '0';
partial_product_23(117) <= '0';
partial_product_23(118) <= '0';
partial_product_23(119) <= '0';
partial_product_23(120) <= '0';
partial_product_23(121) <= '0';
partial_product_23(122) <= '0';
partial_product_23(123) <= '0';
partial_product_23(124) <= '0';
partial_product_23(125) <= '0';
partial_product_23(126) <= '0';
partial_product_23(127) <= '0';
partial_product_23(128) <= '0';
partial_product_23(129) <= '0';
partial_product_23(130) <= '0';
partial_product_23(131) <= '0';
partial_product_23(132) <= '0';
partial_product_23(133) <= '0';
partial_product_23(134) <= '0';
partial_product_23(135) <= '0';
partial_product_23(136) <= '0';
partial_product_23(137) <= '0';
partial_product_23(138) <= '0';
partial_product_23(139) <= '0';
partial_product_23(140) <= '0';
partial_product_23(141) <= '0';
partial_product_23(142) <= '0';
partial_product_23(143) <= '0';
partial_product_23(144) <= '0';
partial_product_23(145) <= '0';
partial_product_23(146) <= '0';
partial_product_23(147) <= '0';
partial_product_23(148) <= '0';
partial_product_23(149) <= '0';
partial_product_23(150) <= '0';
partial_product_23(151) <= '0';
partial_product_23(152) <= '0';
partial_product_23(153) <= '0';
partial_product_23(154) <= '0';
partial_product_23(155) <= '0';
partial_product_23(156) <= '0';
partial_product_23(157) <= '0';
partial_product_23(158) <= '0';
partial_product_23(159) <= '0';
partial_product_23(160) <= '0';
partial_product_23(161) <= '0';
partial_product_23(162) <= '0';
partial_product_23(163) <= '0';
partial_product_23(164) <= '0';
partial_product_23(165) <= '0';
partial_product_23(166) <= '0';
partial_product_23(167) <= '0';
partial_product_23(168) <= '0';
partial_product_23(169) <= '0';
partial_product_23(170) <= '0';
partial_product_23(171) <= '0';
partial_product_23(172) <= '0';
partial_product_23(173) <= '0';
partial_product_23(174) <= '0';
partial_product_23(175) <= '0';
partial_product_23(176) <= '0';
partial_product_23(177) <= '0';
partial_product_23(178) <= '0';
partial_product_23(179) <= '0';
partial_product_23(180) <= '0';
partial_product_23(181) <= '0';
partial_product_23(182) <= '0';
partial_product_23(183) <= '0';
partial_product_23(184) <= '0';
partial_product_23(185) <= '0';
partial_product_23(186) <= '0';
partial_product_23(187) <= '0';
partial_product_23(188) <= '0';
partial_product_23(189) <= '0';
partial_product_23(190) <= '0';
partial_product_23(191) <= '0';
partial_product_23(192) <= '0';
partial_product_23(193) <= '0';
partial_product_23(194) <= '0';
partial_product_23(195) <= '0';
partial_product_23(196) <= '0';
partial_product_23(197) <= '0';
partial_product_23(198) <= '0';
partial_product_23(199) <= '0';
partial_product_23(200) <= '0';
partial_product_23(201) <= '0';
partial_product_23(202) <= '0';
partial_product_23(203) <= '0';
partial_product_23(204) <= '0';
partial_product_23(205) <= '0';
partial_product_23(206) <= '0';
partial_product_23(207) <= '0';
partial_product_23(208) <= '0';
partial_product_23(209) <= '0';
partial_product_23(210) <= '0';
partial_product_23(211) <= '0';
partial_product_23(212) <= '0';
partial_product_23(213) <= '0';
partial_product_23(214) <= '0';
partial_product_23(215) <= '0';
partial_product_23(216) <= '0';
partial_product_23(217) <= '0';
partial_product_23(218) <= '0';
partial_product_23(219) <= '0';
partial_product_23(220) <= '0';
partial_product_23(221) <= '0';
partial_product_23(222) <= '0';
partial_product_23(223) <= '0';
partial_product_23(224) <= '0';
partial_product_23(225) <= '0';
partial_product_23(226) <= '0';
partial_product_23(227) <= '0';
partial_product_23(228) <= '0';
partial_product_23(229) <= '0';
partial_product_23(230) <= '0';
partial_product_23(231) <= '0';
partial_product_23(232) <= '0';
partial_product_23(233) <= '0';
partial_product_23(234) <= '0';
partial_product_23(235) <= '0';
partial_product_23(236) <= '0';
partial_product_23(237) <= '0';
partial_product_23(238) <= temp_mult_86(238);
partial_product_23(239) <= temp_mult_86(239);
partial_product_23(240) <= temp_mult_86(240);
partial_product_23(241) <= temp_mult_86(241);
partial_product_23(242) <= temp_mult_86(242);
partial_product_23(243) <= temp_mult_86(243);
partial_product_23(244) <= temp_mult_86(244);
partial_product_23(245) <= temp_mult_86(245);
partial_product_23(246) <= temp_mult_86(246);
partial_product_23(247) <= temp_mult_86(247);
partial_product_23(248) <= temp_mult_86(248);
partial_product_23(249) <= temp_mult_86(249);
partial_product_23(250) <= temp_mult_86(250);
partial_product_23(251) <= temp_mult_86(251);
partial_product_23(252) <= temp_mult_86(252);
partial_product_23(253) <= temp_mult_86(253);
partial_product_23(254) <= temp_mult_86(254);
partial_product_23(255) <= temp_mult_86(255);
partial_product_23(256) <= temp_mult_86(256);
partial_product_23(257) <= temp_mult_86(257);
partial_product_23(258) <= temp_mult_86(258);
partial_product_23(259) <= temp_mult_86(259);
partial_product_23(260) <= temp_mult_86(260);
partial_product_23(261) <= temp_mult_86(261);
partial_product_23(262) <= temp_mult_86(262);
partial_product_23(263) <= temp_mult_86(263);
partial_product_23(264) <= temp_mult_86(264);
partial_product_23(265) <= temp_mult_86(265);
partial_product_23(266) <= temp_mult_86(266);
partial_product_23(267) <= temp_mult_86(267);
partial_product_23(268) <= temp_mult_86(268);
partial_product_23(269) <= temp_mult_86(269);
partial_product_23(270) <= temp_mult_86(270);
partial_product_23(271) <= temp_mult_86(271);
partial_product_23(272) <= temp_mult_86(272);
partial_product_23(273) <= temp_mult_86(273);
partial_product_23(274) <= temp_mult_86(274);
partial_product_23(275) <= temp_mult_86(275);
partial_product_23(276) <= temp_mult_86(276);
partial_product_23(277) <= temp_mult_86(277);
partial_product_23(278) <= temp_mult_86(278);
partial_product_23(279) <= '0';
partial_product_23(280) <= '0';
partial_product_23(281) <= '0';
partial_product_23(282) <= '0';
partial_product_23(283) <= '0';
partial_product_23(284) <= '0';
partial_product_23(285) <= '0';
partial_product_23(286) <= '0';
partial_product_23(287) <= '0';
partial_product_23(288) <= '0';
partial_product_23(289) <= '0';
partial_product_23(290) <= '0';
partial_product_23(291) <= '0';
partial_product_23(292) <= '0';
partial_product_23(293) <= '0';
partial_product_23(294) <= '0';
partial_product_23(295) <= '0';
partial_product_23(296) <= '0';
partial_product_23(297) <= '0';
partial_product_23(298) <= '0';
partial_product_23(299) <= '0';
partial_product_23(300) <= '0';
partial_product_23(301) <= '0';
partial_product_23(302) <= '0';
partial_product_23(303) <= '0';
partial_product_23(304) <= '0';
partial_product_23(305) <= '0';
partial_product_23(306) <= '0';
partial_product_23(307) <= '0';
partial_product_23(308) <= '0';
partial_product_23(309) <= '0';
partial_product_23(310) <= '0';
partial_product_23(311) <= '0';
partial_product_23(312) <= '0';
partial_product_23(313) <= '0';
partial_product_23(314) <= '0';
partial_product_23(315) <= '0';
partial_product_23(316) <= '0';
partial_product_23(317) <= '0';
partial_product_23(318) <= '0';
partial_product_23(319) <= '0';
partial_product_23(320) <= '0';
partial_product_23(321) <= '0';
partial_product_23(322) <= '0';
partial_product_23(323) <= '0';
partial_product_23(324) <= '0';
partial_product_23(325) <= '0';
partial_product_23(326) <= '0';
partial_product_23(327) <= '0';
partial_product_23(328) <= '0';
partial_product_23(329) <= '0';
partial_product_23(330) <= '0';
partial_product_23(331) <= '0';
partial_product_23(332) <= '0';
partial_product_23(333) <= '0';
partial_product_23(334) <= '0';
partial_product_23(335) <= '0';
partial_product_23(336) <= '0';
partial_product_23(337) <= '0';
partial_product_23(338) <= '0';
partial_product_23(339) <= '0';
partial_product_23(340) <= '0';
partial_product_23(341) <= '0';
partial_product_23(342) <= '0';
partial_product_23(343) <= '0';
partial_product_23(344) <= '0';
partial_product_23(345) <= '0';
partial_product_23(346) <= '0';
partial_product_23(347) <= '0';
partial_product_23(348) <= '0';
partial_product_23(349) <= '0';
partial_product_23(350) <= '0';
partial_product_23(351) <= '0';
partial_product_23(352) <= '0';
partial_product_23(353) <= '0';
partial_product_23(354) <= '0';
partial_product_23(355) <= '0';
partial_product_23(356) <= '0';
partial_product_23(357) <= '0';
partial_product_23(358) <= '0';
partial_product_23(359) <= '0';
partial_product_23(360) <= '0';
partial_product_23(361) <= '0';
partial_product_23(362) <= '0';
partial_product_23(363) <= '0';
partial_product_23(364) <= '0';
partial_product_23(365) <= '0';
partial_product_23(366) <= '0';
partial_product_23(367) <= '0';
partial_product_23(368) <= '0';
partial_product_23(369) <= '0';
partial_product_23(370) <= '0';
partial_product_23(371) <= '0';
partial_product_23(372) <= '0';
partial_product_23(373) <= '0';
partial_product_23(374) <= '0';
partial_product_23(375) <= '0';
partial_product_23(376) <= '0';
partial_product_23(377) <= '0';
partial_product_23(378) <= '0';
partial_product_23(379) <= '0';
partial_product_23(380) <= '0';
partial_product_23(381) <= '0';
partial_product_23(382) <= '0';
partial_product_23(383) <= '0';
partial_product_23(384) <= '0';
partial_product_23(385) <= '0';
partial_product_23(386) <= '0';
partial_product_23(387) <= '0';
partial_product_23(388) <= '0';
partial_product_23(389) <= '0';
partial_product_23(390) <= '0';
partial_product_23(391) <= '0';
partial_product_23(392) <= '0';
partial_product_23(393) <= '0';
partial_product_23(394) <= '0';
partial_product_23(395) <= '0';
partial_product_23(396) <= '0';
partial_product_23(397) <= '0';
partial_product_23(398) <= '0';
partial_product_23(399) <= '0';
partial_product_23(400) <= '0';
partial_product_23(401) <= '0';
partial_product_23(402) <= '0';
partial_product_23(403) <= '0';
partial_product_23(404) <= '0';
partial_product_23(405) <= '0';
partial_product_23(406) <= '0';
partial_product_23(407) <= '0';
partial_product_23(408) <= '0';
partial_product_23(409) <= '0';
partial_product_23(410) <= '0';
partial_product_23(411) <= '0';
partial_product_23(412) <= '0';
partial_product_23(413) <= '0';
partial_product_23(414) <= '0';
partial_product_23(415) <= '0';
partial_product_23(416) <= '0';
partial_product_23(417) <= '0';
partial_product_23(418) <= '0';
partial_product_23(419) <= '0';
partial_product_23(420) <= '0';
partial_product_23(421) <= '0';
partial_product_23(422) <= '0';
partial_product_23(423) <= '0';
partial_product_23(424) <= '0';
partial_product_23(425) <= '0';
partial_product_23(426) <= '0';
partial_product_23(427) <= '0';
partial_product_23(428) <= '0';
partial_product_23(429) <= '0';
partial_product_23(430) <= '0';
partial_product_23(431) <= '0';
partial_product_23(432) <= '0';
partial_product_23(433) <= '0';
partial_product_23(434) <= '0';
partial_product_23(435) <= '0';
partial_product_23(436) <= '0';
partial_product_23(437) <= '0';
partial_product_23(438) <= '0';
partial_product_23(439) <= '0';
partial_product_23(440) <= '0';
partial_product_23(441) <= '0';
partial_product_23(442) <= '0';
partial_product_23(443) <= '0';
partial_product_23(444) <= '0';
partial_product_23(445) <= '0';
partial_product_23(446) <= '0';
partial_product_23(447) <= '0';
partial_product_23(448) <= '0';
partial_product_23(449) <= '0';
partial_product_23(450) <= '0';
partial_product_23(451) <= '0';
partial_product_23(452) <= '0';
partial_product_23(453) <= '0';
partial_product_23(454) <= '0';
partial_product_23(455) <= '0';
partial_product_23(456) <= '0';
partial_product_23(457) <= '0';
partial_product_23(458) <= '0';
partial_product_23(459) <= '0';
partial_product_23(460) <= '0';
partial_product_23(461) <= '0';
partial_product_23(462) <= '0';
partial_product_23(463) <= '0';
partial_product_23(464) <= '0';
partial_product_23(465) <= '0';
partial_product_23(466) <= '0';
partial_product_23(467) <= '0';
partial_product_23(468) <= '0';
partial_product_23(469) <= '0';
partial_product_23(470) <= '0';
partial_product_23(471) <= '0';
partial_product_23(472) <= '0';
partial_product_23(473) <= '0';
partial_product_23(474) <= '0';
partial_product_23(475) <= '0';
partial_product_23(476) <= '0';
partial_product_23(477) <= '0';
partial_product_23(478) <= '0';
partial_product_23(479) <= '0';
partial_product_23(480) <= '0';
partial_product_23(481) <= '0';
partial_product_23(482) <= '0';
partial_product_23(483) <= '0';
partial_product_23(484) <= '0';
partial_product_23(485) <= '0';
partial_product_23(486) <= '0';
partial_product_23(487) <= '0';
partial_product_23(488) <= '0';
partial_product_23(489) <= '0';
partial_product_23(490) <= '0';
partial_product_23(491) <= '0';
partial_product_23(492) <= '0';
partial_product_23(493) <= '0';
partial_product_23(494) <= '0';
partial_product_23(495) <= '0';
partial_product_23(496) <= '0';
partial_product_23(497) <= '0';
partial_product_23(498) <= '0';
partial_product_23(499) <= '0';
partial_product_23(500) <= '0';
partial_product_23(501) <= '0';
partial_product_23(502) <= '0';
partial_product_23(503) <= '0';
partial_product_23(504) <= '0';
partial_product_23(505) <= '0';
partial_product_23(506) <= '0';
partial_product_23(507) <= '0';
partial_product_23(508) <= '0';
partial_product_23(509) <= '0';
partial_product_23(510) <= '0';
partial_product_23(511) <= '0';
partial_product_23(512) <= '0';
partial_product_24(0) <= '0';
partial_product_24(1) <= '0';
partial_product_24(2) <= '0';
partial_product_24(3) <= '0';
partial_product_24(4) <= '0';
partial_product_24(5) <= '0';
partial_product_24(6) <= '0';
partial_product_24(7) <= '0';
partial_product_24(8) <= '0';
partial_product_24(9) <= '0';
partial_product_24(10) <= '0';
partial_product_24(11) <= '0';
partial_product_24(12) <= '0';
partial_product_24(13) <= '0';
partial_product_24(14) <= '0';
partial_product_24(15) <= '0';
partial_product_24(16) <= '0';
partial_product_24(17) <= '0';
partial_product_24(18) <= '0';
partial_product_24(19) <= '0';
partial_product_24(20) <= '0';
partial_product_24(21) <= '0';
partial_product_24(22) <= '0';
partial_product_24(23) <= '0';
partial_product_24(24) <= '0';
partial_product_24(25) <= '0';
partial_product_24(26) <= '0';
partial_product_24(27) <= '0';
partial_product_24(28) <= '0';
partial_product_24(29) <= '0';
partial_product_24(30) <= '0';
partial_product_24(31) <= '0';
partial_product_24(32) <= '0';
partial_product_24(33) <= '0';
partial_product_24(34) <= '0';
partial_product_24(35) <= '0';
partial_product_24(36) <= '0';
partial_product_24(37) <= '0';
partial_product_24(38) <= '0';
partial_product_24(39) <= '0';
partial_product_24(40) <= '0';
partial_product_24(41) <= '0';
partial_product_24(42) <= '0';
partial_product_24(43) <= '0';
partial_product_24(44) <= '0';
partial_product_24(45) <= '0';
partial_product_24(46) <= '0';
partial_product_24(47) <= '0';
partial_product_24(48) <= '0';
partial_product_24(49) <= '0';
partial_product_24(50) <= '0';
partial_product_24(51) <= '0';
partial_product_24(52) <= '0';
partial_product_24(53) <= '0';
partial_product_24(54) <= '0';
partial_product_24(55) <= '0';
partial_product_24(56) <= '0';
partial_product_24(57) <= '0';
partial_product_24(58) <= '0';
partial_product_24(59) <= '0';
partial_product_24(60) <= '0';
partial_product_24(61) <= '0';
partial_product_24(62) <= '0';
partial_product_24(63) <= '0';
partial_product_24(64) <= '0';
partial_product_24(65) <= '0';
partial_product_24(66) <= '0';
partial_product_24(67) <= '0';
partial_product_24(68) <= '0';
partial_product_24(69) <= '0';
partial_product_24(70) <= '0';
partial_product_24(71) <= '0';
partial_product_24(72) <= '0';
partial_product_24(73) <= '0';
partial_product_24(74) <= '0';
partial_product_24(75) <= '0';
partial_product_24(76) <= '0';
partial_product_24(77) <= '0';
partial_product_24(78) <= '0';
partial_product_24(79) <= '0';
partial_product_24(80) <= '0';
partial_product_24(81) <= '0';
partial_product_24(82) <= '0';
partial_product_24(83) <= '0';
partial_product_24(84) <= '0';
partial_product_24(85) <= '0';
partial_product_24(86) <= '0';
partial_product_24(87) <= '0';
partial_product_24(88) <= '0';
partial_product_24(89) <= '0';
partial_product_24(90) <= '0';
partial_product_24(91) <= '0';
partial_product_24(92) <= '0';
partial_product_24(93) <= '0';
partial_product_24(94) <= '0';
partial_product_24(95) <= '0';
partial_product_24(96) <= '0';
partial_product_24(97) <= '0';
partial_product_24(98) <= '0';
partial_product_24(99) <= '0';
partial_product_24(100) <= '0';
partial_product_24(101) <= '0';
partial_product_24(102) <= '0';
partial_product_24(103) <= '0';
partial_product_24(104) <= '0';
partial_product_24(105) <= '0';
partial_product_24(106) <= '0';
partial_product_24(107) <= '0';
partial_product_24(108) <= '0';
partial_product_24(109) <= '0';
partial_product_24(110) <= '0';
partial_product_24(111) <= '0';
partial_product_24(112) <= '0';
partial_product_24(113) <= '0';
partial_product_24(114) <= '0';
partial_product_24(115) <= '0';
partial_product_24(116) <= '0';
partial_product_24(117) <= '0';
partial_product_24(118) <= '0';
partial_product_24(119) <= '0';
partial_product_24(120) <= '0';
partial_product_24(121) <= '0';
partial_product_24(122) <= '0';
partial_product_24(123) <= '0';
partial_product_24(124) <= '0';
partial_product_24(125) <= '0';
partial_product_24(126) <= '0';
partial_product_24(127) <= '0';
partial_product_24(128) <= '0';
partial_product_24(129) <= '0';
partial_product_24(130) <= '0';
partial_product_24(131) <= '0';
partial_product_24(132) <= '0';
partial_product_24(133) <= '0';
partial_product_24(134) <= '0';
partial_product_24(135) <= '0';
partial_product_24(136) <= '0';
partial_product_24(137) <= '0';
partial_product_24(138) <= '0';
partial_product_24(139) <= '0';
partial_product_24(140) <= '0';
partial_product_24(141) <= '0';
partial_product_24(142) <= '0';
partial_product_24(143) <= '0';
partial_product_24(144) <= '0';
partial_product_24(145) <= '0';
partial_product_24(146) <= '0';
partial_product_24(147) <= '0';
partial_product_24(148) <= '0';
partial_product_24(149) <= '0';
partial_product_24(150) <= '0';
partial_product_24(151) <= '0';
partial_product_24(152) <= '0';
partial_product_24(153) <= '0';
partial_product_24(154) <= '0';
partial_product_24(155) <= '0';
partial_product_24(156) <= '0';
partial_product_24(157) <= '0';
partial_product_24(158) <= '0';
partial_product_24(159) <= '0';
partial_product_24(160) <= '0';
partial_product_24(161) <= '0';
partial_product_24(162) <= '0';
partial_product_24(163) <= '0';
partial_product_24(164) <= '0';
partial_product_24(165) <= '0';
partial_product_24(166) <= '0';
partial_product_24(167) <= '0';
partial_product_24(168) <= '0';
partial_product_24(169) <= '0';
partial_product_24(170) <= '0';
partial_product_24(171) <= '0';
partial_product_24(172) <= '0';
partial_product_24(173) <= '0';
partial_product_24(174) <= '0';
partial_product_24(175) <= '0';
partial_product_24(176) <= '0';
partial_product_24(177) <= '0';
partial_product_24(178) <= '0';
partial_product_24(179) <= '0';
partial_product_24(180) <= '0';
partial_product_24(181) <= '0';
partial_product_24(182) <= '0';
partial_product_24(183) <= '0';
partial_product_24(184) <= '0';
partial_product_24(185) <= '0';
partial_product_24(186) <= '0';
partial_product_24(187) <= '0';
partial_product_24(188) <= '0';
partial_product_24(189) <= '0';
partial_product_24(190) <= '0';
partial_product_24(191) <= '0';
partial_product_24(192) <= '0';
partial_product_24(193) <= '0';
partial_product_24(194) <= '0';
partial_product_24(195) <= '0';
partial_product_24(196) <= '0';
partial_product_24(197) <= '0';
partial_product_24(198) <= '0';
partial_product_24(199) <= '0';
partial_product_24(200) <= '0';
partial_product_24(201) <= '0';
partial_product_24(202) <= '0';
partial_product_24(203) <= '0';
partial_product_24(204) <= '0';
partial_product_24(205) <= '0';
partial_product_24(206) <= '0';
partial_product_24(207) <= '0';
partial_product_24(208) <= '0';
partial_product_24(209) <= '0';
partial_product_24(210) <= '0';
partial_product_24(211) <= '0';
partial_product_24(212) <= '0';
partial_product_24(213) <= '0';
partial_product_24(214) <= '0';
partial_product_24(215) <= '0';
partial_product_24(216) <= '0';
partial_product_24(217) <= '0';
partial_product_24(218) <= '0';
partial_product_24(219) <= '0';
partial_product_24(220) <= '0';
partial_product_24(221) <= '0';
partial_product_24(222) <= '0';
partial_product_24(223) <= '0';
partial_product_24(224) <= '0';
partial_product_24(225) <= '0';
partial_product_24(226) <= '0';
partial_product_24(227) <= '0';
partial_product_24(228) <= '0';
partial_product_24(229) <= '0';
partial_product_24(230) <= '0';
partial_product_24(231) <= '0';
partial_product_24(232) <= '0';
partial_product_24(233) <= '0';
partial_product_24(234) <= '0';
partial_product_24(235) <= '0';
partial_product_24(236) <= '0';
partial_product_24(237) <= '0';
partial_product_24(238) <= '0';
partial_product_24(239) <= '0';
partial_product_24(240) <= temp_mult_160(240);
partial_product_24(241) <= temp_mult_160(241);
partial_product_24(242) <= temp_mult_160(242);
partial_product_24(243) <= temp_mult_160(243);
partial_product_24(244) <= temp_mult_160(244);
partial_product_24(245) <= temp_mult_160(245);
partial_product_24(246) <= temp_mult_160(246);
partial_product_24(247) <= temp_mult_160(247);
partial_product_24(248) <= temp_mult_160(248);
partial_product_24(249) <= temp_mult_160(249);
partial_product_24(250) <= temp_mult_160(250);
partial_product_24(251) <= temp_mult_160(251);
partial_product_24(252) <= temp_mult_160(252);
partial_product_24(253) <= temp_mult_160(253);
partial_product_24(254) <= temp_mult_160(254);
partial_product_24(255) <= temp_mult_160(255);
partial_product_24(256) <= temp_mult_160(256);
partial_product_24(257) <= temp_mult_160(257);
partial_product_24(258) <= temp_mult_160(258);
partial_product_24(259) <= temp_mult_160(259);
partial_product_24(260) <= temp_mult_160(260);
partial_product_24(261) <= temp_mult_160(261);
partial_product_24(262) <= temp_mult_160(262);
partial_product_24(263) <= temp_mult_160(263);
partial_product_24(264) <= temp_mult_160(264);
partial_product_24(265) <= temp_mult_160(265);
partial_product_24(266) <= temp_mult_160(266);
partial_product_24(267) <= temp_mult_160(267);
partial_product_24(268) <= temp_mult_160(268);
partial_product_24(269) <= temp_mult_160(269);
partial_product_24(270) <= temp_mult_160(270);
partial_product_24(271) <= temp_mult_160(271);
partial_product_24(272) <= '0';
partial_product_24(273) <= '0';
partial_product_24(274) <= '0';
partial_product_24(275) <= '0';
partial_product_24(276) <= '0';
partial_product_24(277) <= '0';
partial_product_24(278) <= '0';
partial_product_24(279) <= '0';
partial_product_24(280) <= '0';
partial_product_24(281) <= '0';
partial_product_24(282) <= '0';
partial_product_24(283) <= '0';
partial_product_24(284) <= '0';
partial_product_24(285) <= '0';
partial_product_24(286) <= '0';
partial_product_24(287) <= '0';
partial_product_24(288) <= '0';
partial_product_24(289) <= '0';
partial_product_24(290) <= '0';
partial_product_24(291) <= '0';
partial_product_24(292) <= '0';
partial_product_24(293) <= '0';
partial_product_24(294) <= '0';
partial_product_24(295) <= '0';
partial_product_24(296) <= '0';
partial_product_24(297) <= '0';
partial_product_24(298) <= '0';
partial_product_24(299) <= '0';
partial_product_24(300) <= '0';
partial_product_24(301) <= '0';
partial_product_24(302) <= '0';
partial_product_24(303) <= '0';
partial_product_24(304) <= '0';
partial_product_24(305) <= '0';
partial_product_24(306) <= '0';
partial_product_24(307) <= '0';
partial_product_24(308) <= '0';
partial_product_24(309) <= '0';
partial_product_24(310) <= '0';
partial_product_24(311) <= '0';
partial_product_24(312) <= '0';
partial_product_24(313) <= '0';
partial_product_24(314) <= '0';
partial_product_24(315) <= '0';
partial_product_24(316) <= '0';
partial_product_24(317) <= '0';
partial_product_24(318) <= '0';
partial_product_24(319) <= '0';
partial_product_24(320) <= '0';
partial_product_24(321) <= '0';
partial_product_24(322) <= '0';
partial_product_24(323) <= '0';
partial_product_24(324) <= '0';
partial_product_24(325) <= '0';
partial_product_24(326) <= '0';
partial_product_24(327) <= '0';
partial_product_24(328) <= '0';
partial_product_24(329) <= '0';
partial_product_24(330) <= '0';
partial_product_24(331) <= '0';
partial_product_24(332) <= '0';
partial_product_24(333) <= '0';
partial_product_24(334) <= '0';
partial_product_24(335) <= '0';
partial_product_24(336) <= '0';
partial_product_24(337) <= '0';
partial_product_24(338) <= '0';
partial_product_24(339) <= '0';
partial_product_24(340) <= '0';
partial_product_24(341) <= '0';
partial_product_24(342) <= '0';
partial_product_24(343) <= '0';
partial_product_24(344) <= '0';
partial_product_24(345) <= '0';
partial_product_24(346) <= '0';
partial_product_24(347) <= '0';
partial_product_24(348) <= '0';
partial_product_24(349) <= '0';
partial_product_24(350) <= '0';
partial_product_24(351) <= '0';
partial_product_24(352) <= '0';
partial_product_24(353) <= '0';
partial_product_24(354) <= '0';
partial_product_24(355) <= '0';
partial_product_24(356) <= '0';
partial_product_24(357) <= '0';
partial_product_24(358) <= '0';
partial_product_24(359) <= '0';
partial_product_24(360) <= '0';
partial_product_24(361) <= '0';
partial_product_24(362) <= '0';
partial_product_24(363) <= '0';
partial_product_24(364) <= '0';
partial_product_24(365) <= '0';
partial_product_24(366) <= '0';
partial_product_24(367) <= '0';
partial_product_24(368) <= '0';
partial_product_24(369) <= '0';
partial_product_24(370) <= '0';
partial_product_24(371) <= '0';
partial_product_24(372) <= '0';
partial_product_24(373) <= '0';
partial_product_24(374) <= '0';
partial_product_24(375) <= '0';
partial_product_24(376) <= '0';
partial_product_24(377) <= '0';
partial_product_24(378) <= '0';
partial_product_24(379) <= '0';
partial_product_24(380) <= '0';
partial_product_24(381) <= '0';
partial_product_24(382) <= '0';
partial_product_24(383) <= '0';
partial_product_24(384) <= '0';
partial_product_24(385) <= '0';
partial_product_24(386) <= '0';
partial_product_24(387) <= '0';
partial_product_24(388) <= '0';
partial_product_24(389) <= '0';
partial_product_24(390) <= '0';
partial_product_24(391) <= '0';
partial_product_24(392) <= '0';
partial_product_24(393) <= '0';
partial_product_24(394) <= '0';
partial_product_24(395) <= '0';
partial_product_24(396) <= '0';
partial_product_24(397) <= '0';
partial_product_24(398) <= '0';
partial_product_24(399) <= '0';
partial_product_24(400) <= '0';
partial_product_24(401) <= '0';
partial_product_24(402) <= '0';
partial_product_24(403) <= '0';
partial_product_24(404) <= '0';
partial_product_24(405) <= '0';
partial_product_24(406) <= '0';
partial_product_24(407) <= '0';
partial_product_24(408) <= '0';
partial_product_24(409) <= '0';
partial_product_24(410) <= '0';
partial_product_24(411) <= '0';
partial_product_24(412) <= '0';
partial_product_24(413) <= '0';
partial_product_24(414) <= '0';
partial_product_24(415) <= '0';
partial_product_24(416) <= '0';
partial_product_24(417) <= '0';
partial_product_24(418) <= '0';
partial_product_24(419) <= '0';
partial_product_24(420) <= '0';
partial_product_24(421) <= '0';
partial_product_24(422) <= '0';
partial_product_24(423) <= '0';
partial_product_24(424) <= '0';
partial_product_24(425) <= '0';
partial_product_24(426) <= '0';
partial_product_24(427) <= '0';
partial_product_24(428) <= '0';
partial_product_24(429) <= '0';
partial_product_24(430) <= '0';
partial_product_24(431) <= '0';
partial_product_24(432) <= '0';
partial_product_24(433) <= '0';
partial_product_24(434) <= '0';
partial_product_24(435) <= '0';
partial_product_24(436) <= '0';
partial_product_24(437) <= '0';
partial_product_24(438) <= '0';
partial_product_24(439) <= '0';
partial_product_24(440) <= '0';
partial_product_24(441) <= '0';
partial_product_24(442) <= '0';
partial_product_24(443) <= '0';
partial_product_24(444) <= '0';
partial_product_24(445) <= '0';
partial_product_24(446) <= '0';
partial_product_24(447) <= '0';
partial_product_24(448) <= '0';
partial_product_24(449) <= '0';
partial_product_24(450) <= '0';
partial_product_24(451) <= '0';
partial_product_24(452) <= '0';
partial_product_24(453) <= '0';
partial_product_24(454) <= '0';
partial_product_24(455) <= '0';
partial_product_24(456) <= '0';
partial_product_24(457) <= '0';
partial_product_24(458) <= '0';
partial_product_24(459) <= '0';
partial_product_24(460) <= '0';
partial_product_24(461) <= '0';
partial_product_24(462) <= '0';
partial_product_24(463) <= '0';
partial_product_24(464) <= '0';
partial_product_24(465) <= '0';
partial_product_24(466) <= '0';
partial_product_24(467) <= '0';
partial_product_24(468) <= '0';
partial_product_24(469) <= '0';
partial_product_24(470) <= '0';
partial_product_24(471) <= '0';
partial_product_24(472) <= '0';
partial_product_24(473) <= '0';
partial_product_24(474) <= '0';
partial_product_24(475) <= '0';
partial_product_24(476) <= '0';
partial_product_24(477) <= '0';
partial_product_24(478) <= '0';
partial_product_24(479) <= '0';
partial_product_24(480) <= '0';
partial_product_24(481) <= '0';
partial_product_24(482) <= '0';
partial_product_24(483) <= '0';
partial_product_24(484) <= '0';
partial_product_24(485) <= '0';
partial_product_24(486) <= '0';
partial_product_24(487) <= '0';
partial_product_24(488) <= '0';
partial_product_24(489) <= '0';
partial_product_24(490) <= '0';
partial_product_24(491) <= '0';
partial_product_24(492) <= '0';
partial_product_24(493) <= '0';
partial_product_24(494) <= '0';
partial_product_24(495) <= '0';
partial_product_24(496) <= '0';
partial_product_24(497) <= '0';
partial_product_24(498) <= '0';
partial_product_24(499) <= '0';
partial_product_24(500) <= '0';
partial_product_24(501) <= '0';
partial_product_24(502) <= '0';
partial_product_24(503) <= '0';
partial_product_24(504) <= '0';
partial_product_24(505) <= '0';
partial_product_24(506) <= '0';
partial_product_24(507) <= '0';
partial_product_24(508) <= '0';
partial_product_24(509) <= '0';
partial_product_24(510) <= '0';
partial_product_24(511) <= '0';
partial_product_24(512) <= '0';
partial_product_25(0) <= '0';
partial_product_25(1) <= '0';
partial_product_25(2) <= '0';
partial_product_25(3) <= '0';
partial_product_25(4) <= '0';
partial_product_25(5) <= '0';
partial_product_25(6) <= '0';
partial_product_25(7) <= '0';
partial_product_25(8) <= '0';
partial_product_25(9) <= '0';
partial_product_25(10) <= '0';
partial_product_25(11) <= '0';
partial_product_25(12) <= '0';
partial_product_25(13) <= '0';
partial_product_25(14) <= '0';
partial_product_25(15) <= '0';
partial_product_25(16) <= '0';
partial_product_25(17) <= '0';
partial_product_25(18) <= '0';
partial_product_25(19) <= '0';
partial_product_25(20) <= '0';
partial_product_25(21) <= '0';
partial_product_25(22) <= '0';
partial_product_25(23) <= '0';
partial_product_25(24) <= '0';
partial_product_25(25) <= '0';
partial_product_25(26) <= '0';
partial_product_25(27) <= '0';
partial_product_25(28) <= '0';
partial_product_25(29) <= '0';
partial_product_25(30) <= '0';
partial_product_25(31) <= '0';
partial_product_25(32) <= '0';
partial_product_25(33) <= '0';
partial_product_25(34) <= '0';
partial_product_25(35) <= '0';
partial_product_25(36) <= '0';
partial_product_25(37) <= '0';
partial_product_25(38) <= '0';
partial_product_25(39) <= '0';
partial_product_25(40) <= '0';
partial_product_25(41) <= '0';
partial_product_25(42) <= '0';
partial_product_25(43) <= '0';
partial_product_25(44) <= '0';
partial_product_25(45) <= '0';
partial_product_25(46) <= '0';
partial_product_25(47) <= '0';
partial_product_25(48) <= '0';
partial_product_25(49) <= '0';
partial_product_25(50) <= '0';
partial_product_25(51) <= '0';
partial_product_25(52) <= '0';
partial_product_25(53) <= '0';
partial_product_25(54) <= '0';
partial_product_25(55) <= '0';
partial_product_25(56) <= '0';
partial_product_25(57) <= '0';
partial_product_25(58) <= '0';
partial_product_25(59) <= '0';
partial_product_25(60) <= '0';
partial_product_25(61) <= '0';
partial_product_25(62) <= '0';
partial_product_25(63) <= '0';
partial_product_25(64) <= '0';
partial_product_25(65) <= '0';
partial_product_25(66) <= '0';
partial_product_25(67) <= '0';
partial_product_25(68) <= '0';
partial_product_25(69) <= '0';
partial_product_25(70) <= '0';
partial_product_25(71) <= '0';
partial_product_25(72) <= '0';
partial_product_25(73) <= '0';
partial_product_25(74) <= '0';
partial_product_25(75) <= '0';
partial_product_25(76) <= '0';
partial_product_25(77) <= '0';
partial_product_25(78) <= '0';
partial_product_25(79) <= '0';
partial_product_25(80) <= '0';
partial_product_25(81) <= '0';
partial_product_25(82) <= '0';
partial_product_25(83) <= '0';
partial_product_25(84) <= '0';
partial_product_25(85) <= '0';
partial_product_25(86) <= '0';
partial_product_25(87) <= '0';
partial_product_25(88) <= '0';
partial_product_25(89) <= '0';
partial_product_25(90) <= '0';
partial_product_25(91) <= '0';
partial_product_25(92) <= '0';
partial_product_25(93) <= '0';
partial_product_25(94) <= '0';
partial_product_25(95) <= '0';
partial_product_25(96) <= '0';
partial_product_25(97) <= '0';
partial_product_25(98) <= '0';
partial_product_25(99) <= '0';
partial_product_25(100) <= '0';
partial_product_25(101) <= '0';
partial_product_25(102) <= '0';
partial_product_25(103) <= '0';
partial_product_25(104) <= '0';
partial_product_25(105) <= '0';
partial_product_25(106) <= '0';
partial_product_25(107) <= '0';
partial_product_25(108) <= '0';
partial_product_25(109) <= '0';
partial_product_25(110) <= '0';
partial_product_25(111) <= '0';
partial_product_25(112) <= '0';
partial_product_25(113) <= '0';
partial_product_25(114) <= '0';
partial_product_25(115) <= '0';
partial_product_25(116) <= '0';
partial_product_25(117) <= '0';
partial_product_25(118) <= '0';
partial_product_25(119) <= '0';
partial_product_25(120) <= '0';
partial_product_25(121) <= '0';
partial_product_25(122) <= '0';
partial_product_25(123) <= '0';
partial_product_25(124) <= '0';
partial_product_25(125) <= '0';
partial_product_25(126) <= '0';
partial_product_25(127) <= '0';
partial_product_25(128) <= '0';
partial_product_25(129) <= '0';
partial_product_25(130) <= '0';
partial_product_25(131) <= '0';
partial_product_25(132) <= '0';
partial_product_25(133) <= '0';
partial_product_25(134) <= '0';
partial_product_25(135) <= '0';
partial_product_25(136) <= '0';
partial_product_25(137) <= '0';
partial_product_25(138) <= '0';
partial_product_25(139) <= '0';
partial_product_25(140) <= '0';
partial_product_25(141) <= '0';
partial_product_25(142) <= '0';
partial_product_25(143) <= '0';
partial_product_25(144) <= '0';
partial_product_25(145) <= '0';
partial_product_25(146) <= '0';
partial_product_25(147) <= '0';
partial_product_25(148) <= '0';
partial_product_25(149) <= '0';
partial_product_25(150) <= '0';
partial_product_25(151) <= '0';
partial_product_25(152) <= '0';
partial_product_25(153) <= '0';
partial_product_25(154) <= '0';
partial_product_25(155) <= '0';
partial_product_25(156) <= '0';
partial_product_25(157) <= '0';
partial_product_25(158) <= '0';
partial_product_25(159) <= '0';
partial_product_25(160) <= '0';
partial_product_25(161) <= '0';
partial_product_25(162) <= '0';
partial_product_25(163) <= '0';
partial_product_25(164) <= '0';
partial_product_25(165) <= '0';
partial_product_25(166) <= '0';
partial_product_25(167) <= '0';
partial_product_25(168) <= '0';
partial_product_25(169) <= '0';
partial_product_25(170) <= '0';
partial_product_25(171) <= '0';
partial_product_25(172) <= '0';
partial_product_25(173) <= '0';
partial_product_25(174) <= '0';
partial_product_25(175) <= '0';
partial_product_25(176) <= '0';
partial_product_25(177) <= '0';
partial_product_25(178) <= '0';
partial_product_25(179) <= '0';
partial_product_25(180) <= '0';
partial_product_25(181) <= '0';
partial_product_25(182) <= '0';
partial_product_25(183) <= '0';
partial_product_25(184) <= '0';
partial_product_25(185) <= '0';
partial_product_25(186) <= '0';
partial_product_25(187) <= '0';
partial_product_25(188) <= '0';
partial_product_25(189) <= '0';
partial_product_25(190) <= '0';
partial_product_25(191) <= '0';
partial_product_25(192) <= '0';
partial_product_25(193) <= '0';
partial_product_25(194) <= '0';
partial_product_25(195) <= '0';
partial_product_25(196) <= '0';
partial_product_25(197) <= '0';
partial_product_25(198) <= '0';
partial_product_25(199) <= '0';
partial_product_25(200) <= '0';
partial_product_25(201) <= '0';
partial_product_25(202) <= '0';
partial_product_25(203) <= '0';
partial_product_25(204) <= '0';
partial_product_25(205) <= '0';
partial_product_25(206) <= '0';
partial_product_25(207) <= '0';
partial_product_25(208) <= '0';
partial_product_25(209) <= '0';
partial_product_25(210) <= '0';
partial_product_25(211) <= '0';
partial_product_25(212) <= '0';
partial_product_25(213) <= '0';
partial_product_25(214) <= '0';
partial_product_25(215) <= '0';
partial_product_25(216) <= '0';
partial_product_25(217) <= '0';
partial_product_25(218) <= '0';
partial_product_25(219) <= '0';
partial_product_25(220) <= '0';
partial_product_25(221) <= '0';
partial_product_25(222) <= '0';
partial_product_25(223) <= '0';
partial_product_25(224) <= '0';
partial_product_25(225) <= '0';
partial_product_25(226) <= '0';
partial_product_25(227) <= '0';
partial_product_25(228) <= '0';
partial_product_25(229) <= '0';
partial_product_25(230) <= '0';
partial_product_25(231) <= '0';
partial_product_25(232) <= '0';
partial_product_25(233) <= '0';
partial_product_25(234) <= '0';
partial_product_25(235) <= '0';
partial_product_25(236) <= '0';
partial_product_25(237) <= '0';
partial_product_25(238) <= '0';
partial_product_25(239) <= '0';
partial_product_25(240) <= '0';
partial_product_25(241) <= '0';
partial_product_25(242) <= '0';
partial_product_25(243) <= '0';
partial_product_25(244) <= '0';
partial_product_25(245) <= '0';
partial_product_25(246) <= '0';
partial_product_25(247) <= '0';
partial_product_25(248) <= '0';
partial_product_25(249) <= '0';
partial_product_25(250) <= '0';
partial_product_25(251) <= '0';
partial_product_25(252) <= '0';
partial_product_25(253) <= '0';
partial_product_25(254) <= '0';
partial_product_25(255) <= temp_mult_87(255);
partial_product_25(256) <= temp_mult_87(256);
partial_product_25(257) <= temp_mult_87(257);
partial_product_25(258) <= temp_mult_87(258);
partial_product_25(259) <= temp_mult_87(259);
partial_product_25(260) <= temp_mult_87(260);
partial_product_25(261) <= temp_mult_87(261);
partial_product_25(262) <= temp_mult_87(262);
partial_product_25(263) <= temp_mult_87(263);
partial_product_25(264) <= temp_mult_87(264);
partial_product_25(265) <= temp_mult_87(265);
partial_product_25(266) <= temp_mult_87(266);
partial_product_25(267) <= temp_mult_87(267);
partial_product_25(268) <= temp_mult_87(268);
partial_product_25(269) <= temp_mult_87(269);
partial_product_25(270) <= temp_mult_87(270);
partial_product_25(271) <= temp_mult_87(271);
partial_product_25(272) <= temp_mult_87(272);
partial_product_25(273) <= temp_mult_87(273);
partial_product_25(274) <= temp_mult_87(274);
partial_product_25(275) <= temp_mult_87(275);
partial_product_25(276) <= temp_mult_87(276);
partial_product_25(277) <= temp_mult_87(277);
partial_product_25(278) <= temp_mult_87(278);
partial_product_25(279) <= temp_mult_87(279);
partial_product_25(280) <= temp_mult_87(280);
partial_product_25(281) <= temp_mult_87(281);
partial_product_25(282) <= temp_mult_87(282);
partial_product_25(283) <= temp_mult_87(283);
partial_product_25(284) <= temp_mult_87(284);
partial_product_25(285) <= temp_mult_87(285);
partial_product_25(286) <= temp_mult_87(286);
partial_product_25(287) <= temp_mult_87(287);
partial_product_25(288) <= temp_mult_87(288);
partial_product_25(289) <= temp_mult_87(289);
partial_product_25(290) <= temp_mult_87(290);
partial_product_25(291) <= temp_mult_87(291);
partial_product_25(292) <= temp_mult_87(292);
partial_product_25(293) <= temp_mult_87(293);
partial_product_25(294) <= temp_mult_87(294);
partial_product_25(295) <= temp_mult_87(295);
partial_product_25(296) <= '0';
partial_product_25(297) <= '0';
partial_product_25(298) <= '0';
partial_product_25(299) <= '0';
partial_product_25(300) <= '0';
partial_product_25(301) <= '0';
partial_product_25(302) <= '0';
partial_product_25(303) <= '0';
partial_product_25(304) <= '0';
partial_product_25(305) <= '0';
partial_product_25(306) <= '0';
partial_product_25(307) <= '0';
partial_product_25(308) <= '0';
partial_product_25(309) <= '0';
partial_product_25(310) <= '0';
partial_product_25(311) <= '0';
partial_product_25(312) <= '0';
partial_product_25(313) <= '0';
partial_product_25(314) <= '0';
partial_product_25(315) <= '0';
partial_product_25(316) <= '0';
partial_product_25(317) <= '0';
partial_product_25(318) <= '0';
partial_product_25(319) <= '0';
partial_product_25(320) <= '0';
partial_product_25(321) <= '0';
partial_product_25(322) <= '0';
partial_product_25(323) <= '0';
partial_product_25(324) <= '0';
partial_product_25(325) <= '0';
partial_product_25(326) <= '0';
partial_product_25(327) <= '0';
partial_product_25(328) <= '0';
partial_product_25(329) <= '0';
partial_product_25(330) <= '0';
partial_product_25(331) <= '0';
partial_product_25(332) <= '0';
partial_product_25(333) <= '0';
partial_product_25(334) <= '0';
partial_product_25(335) <= '0';
partial_product_25(336) <= '0';
partial_product_25(337) <= '0';
partial_product_25(338) <= '0';
partial_product_25(339) <= '0';
partial_product_25(340) <= '0';
partial_product_25(341) <= '0';
partial_product_25(342) <= '0';
partial_product_25(343) <= '0';
partial_product_25(344) <= '0';
partial_product_25(345) <= '0';
partial_product_25(346) <= '0';
partial_product_25(347) <= '0';
partial_product_25(348) <= '0';
partial_product_25(349) <= '0';
partial_product_25(350) <= '0';
partial_product_25(351) <= '0';
partial_product_25(352) <= '0';
partial_product_25(353) <= '0';
partial_product_25(354) <= '0';
partial_product_25(355) <= '0';
partial_product_25(356) <= '0';
partial_product_25(357) <= '0';
partial_product_25(358) <= '0';
partial_product_25(359) <= '0';
partial_product_25(360) <= '0';
partial_product_25(361) <= '0';
partial_product_25(362) <= '0';
partial_product_25(363) <= '0';
partial_product_25(364) <= '0';
partial_product_25(365) <= '0';
partial_product_25(366) <= '0';
partial_product_25(367) <= '0';
partial_product_25(368) <= '0';
partial_product_25(369) <= '0';
partial_product_25(370) <= '0';
partial_product_25(371) <= '0';
partial_product_25(372) <= '0';
partial_product_25(373) <= '0';
partial_product_25(374) <= '0';
partial_product_25(375) <= '0';
partial_product_25(376) <= '0';
partial_product_25(377) <= '0';
partial_product_25(378) <= '0';
partial_product_25(379) <= '0';
partial_product_25(380) <= '0';
partial_product_25(381) <= '0';
partial_product_25(382) <= '0';
partial_product_25(383) <= '0';
partial_product_25(384) <= '0';
partial_product_25(385) <= '0';
partial_product_25(386) <= '0';
partial_product_25(387) <= '0';
partial_product_25(388) <= '0';
partial_product_25(389) <= '0';
partial_product_25(390) <= '0';
partial_product_25(391) <= '0';
partial_product_25(392) <= '0';
partial_product_25(393) <= '0';
partial_product_25(394) <= '0';
partial_product_25(395) <= '0';
partial_product_25(396) <= '0';
partial_product_25(397) <= '0';
partial_product_25(398) <= '0';
partial_product_25(399) <= '0';
partial_product_25(400) <= '0';
partial_product_25(401) <= '0';
partial_product_25(402) <= '0';
partial_product_25(403) <= '0';
partial_product_25(404) <= '0';
partial_product_25(405) <= '0';
partial_product_25(406) <= '0';
partial_product_25(407) <= '0';
partial_product_25(408) <= '0';
partial_product_25(409) <= '0';
partial_product_25(410) <= '0';
partial_product_25(411) <= '0';
partial_product_25(412) <= '0';
partial_product_25(413) <= '0';
partial_product_25(414) <= '0';
partial_product_25(415) <= '0';
partial_product_25(416) <= '0';
partial_product_25(417) <= '0';
partial_product_25(418) <= '0';
partial_product_25(419) <= '0';
partial_product_25(420) <= '0';
partial_product_25(421) <= '0';
partial_product_25(422) <= '0';
partial_product_25(423) <= '0';
partial_product_25(424) <= '0';
partial_product_25(425) <= '0';
partial_product_25(426) <= '0';
partial_product_25(427) <= '0';
partial_product_25(428) <= '0';
partial_product_25(429) <= '0';
partial_product_25(430) <= '0';
partial_product_25(431) <= '0';
partial_product_25(432) <= '0';
partial_product_25(433) <= '0';
partial_product_25(434) <= '0';
partial_product_25(435) <= '0';
partial_product_25(436) <= '0';
partial_product_25(437) <= '0';
partial_product_25(438) <= '0';
partial_product_25(439) <= '0';
partial_product_25(440) <= '0';
partial_product_25(441) <= '0';
partial_product_25(442) <= '0';
partial_product_25(443) <= '0';
partial_product_25(444) <= '0';
partial_product_25(445) <= '0';
partial_product_25(446) <= '0';
partial_product_25(447) <= '0';
partial_product_25(448) <= '0';
partial_product_25(449) <= '0';
partial_product_25(450) <= '0';
partial_product_25(451) <= '0';
partial_product_25(452) <= '0';
partial_product_25(453) <= '0';
partial_product_25(454) <= '0';
partial_product_25(455) <= '0';
partial_product_25(456) <= '0';
partial_product_25(457) <= '0';
partial_product_25(458) <= '0';
partial_product_25(459) <= '0';
partial_product_25(460) <= '0';
partial_product_25(461) <= '0';
partial_product_25(462) <= '0';
partial_product_25(463) <= '0';
partial_product_25(464) <= '0';
partial_product_25(465) <= '0';
partial_product_25(466) <= '0';
partial_product_25(467) <= '0';
partial_product_25(468) <= '0';
partial_product_25(469) <= '0';
partial_product_25(470) <= '0';
partial_product_25(471) <= '0';
partial_product_25(472) <= '0';
partial_product_25(473) <= '0';
partial_product_25(474) <= '0';
partial_product_25(475) <= '0';
partial_product_25(476) <= '0';
partial_product_25(477) <= '0';
partial_product_25(478) <= '0';
partial_product_25(479) <= '0';
partial_product_25(480) <= '0';
partial_product_25(481) <= '0';
partial_product_25(482) <= '0';
partial_product_25(483) <= '0';
partial_product_25(484) <= '0';
partial_product_25(485) <= '0';
partial_product_25(486) <= '0';
partial_product_25(487) <= '0';
partial_product_25(488) <= '0';
partial_product_25(489) <= '0';
partial_product_25(490) <= '0';
partial_product_25(491) <= '0';
partial_product_25(492) <= '0';
partial_product_25(493) <= '0';
partial_product_25(494) <= '0';
partial_product_25(495) <= '0';
partial_product_25(496) <= '0';
partial_product_25(497) <= '0';
partial_product_25(498) <= '0';
partial_product_25(499) <= '0';
partial_product_25(500) <= '0';
partial_product_25(501) <= '0';
partial_product_25(502) <= '0';
partial_product_25(503) <= '0';
partial_product_25(504) <= '0';
partial_product_25(505) <= '0';
partial_product_25(506) <= '0';
partial_product_25(507) <= '0';
partial_product_25(508) <= '0';
partial_product_25(509) <= '0';
partial_product_25(510) <= '0';
partial_product_25(511) <= '0';
partial_product_25(512) <= '0';

partial_product_26(255 downto 0) <= (others => '0');
partial_product_26(513 downto 256) <= temp_mult_161;

partial_product_27(255 downto 0) <= (others => '0');
partial_product_27(513 downto 256) <= temp_mult_162;

process(clk)
begin
    if(rising_edge(clk)) then
        temp_o1 <= (signed(partial_product_0) + signed(partial_product_1) + signed(partial_product_2) + signed(partial_product_3) + signed(partial_product_4) + signed(partial_product_5) + signed(partial_product_6) + signed(partial_product_7) + signed(partial_product_8) + signed(partial_product_9) + signed(partial_product_10) + signed(partial_product_11) + signed(partial_product_12) + signed(partial_product_13) + signed(partial_product_14) + signed(partial_product_15) + signed(partial_product_16) + signed(partial_product_17) + signed(partial_product_18) + signed(partial_product_19) + signed(partial_product_20) + signed(partial_product_21) + signed(partial_product_22) + signed(partial_product_23) + signed(partial_product_24) + signed(partial_product_25) - signed(partial_product_26) - signed(partial_product_27));
        temp_o2 <= temp_o1;
        temp_o3 <= temp_o2;
        temp_o4 <= temp_o3;
        temp_o5 <= temp_o4;
        o <= std_logic_vector(temp_o5);
    end if;
end process;

end tiled_behavioral_v1;

















































architecture tiled_behavioral_v2 of pipeline_signed_base_multiplier_257 is

component adder_compressor_30_5
    Generic(
        total_size : integer
    );
    Port (
        a1 : in std_logic_vector((total_size - 1) downto 0);
        a2 : in std_logic_vector((total_size - 1) downto 0);
        a3 : in std_logic_vector((total_size - 1) downto 0);
        a4 : in std_logic_vector((total_size - 1) downto 0);
        a5 : in std_logic_vector((total_size - 1) downto 0);
        a6 : in std_logic_vector((total_size - 1) downto 0);
        a7 : in std_logic_vector((total_size - 1) downto 0);
        a8 : in std_logic_vector((total_size - 1) downto 0);
        a9 : in std_logic_vector((total_size - 1) downto 0);
        a10 : in std_logic_vector((total_size - 1) downto 0);
        a11 : in std_logic_vector((total_size - 1) downto 0);
        a12 : in std_logic_vector((total_size - 1) downto 0);
        a13 : in std_logic_vector((total_size - 1) downto 0);
        a14 : in std_logic_vector((total_size - 1) downto 0);
        a15 : in std_logic_vector((total_size - 1) downto 0);
        a16 : in std_logic_vector((total_size - 1) downto 0);
        a17 : in std_logic_vector((total_size - 1) downto 0);
        a18 : in std_logic_vector((total_size - 1) downto 0);
        a19 : in std_logic_vector((total_size - 1) downto 0);
        a20 : in std_logic_vector((total_size - 1) downto 0);
        a21 : in std_logic_vector((total_size - 1) downto 0);
        a22 : in std_logic_vector((total_size - 1) downto 0);
        a23 : in std_logic_vector((total_size - 1) downto 0);
        a24 : in std_logic_vector((total_size - 1) downto 0);
        a25 : in std_logic_vector((total_size - 1) downto 0);
        a26 : in std_logic_vector((total_size - 1) downto 0);
        a27 : in std_logic_vector((total_size - 1) downto 0);
        a28 : in std_logic_vector((total_size - 1) downto 0);
        a29 : in std_logic_vector((total_size - 1) downto 0);
        a30 : in std_logic_vector((total_size - 1) downto 0);
        c1 : out std_logic_vector((total_size) downto 0);
        c2 : out std_logic_vector((total_size+1) downto 0);
        c3 : out std_logic_vector((total_size+2) downto 0);
        c4 : out std_logic_vector((total_size+3) downto 0);
        s : out std_logic_vector((total_size - 1) downto 0)
    );
end component;

component adder_compressor_5_3
    Generic(
        total_size : integer
    );
    Port (
        a1 : in std_logic_vector((total_size - 1) downto 0);
        a2 : in std_logic_vector((total_size - 1) downto 0);
        a3 : in std_logic_vector((total_size - 1) downto 0);
        a4 : in std_logic_vector((total_size - 1) downto 0);
        a5 : in std_logic_vector((total_size - 1) downto 0);
        c1 : out std_logic_vector((total_size) downto 0);
        c2 : out std_logic_vector((total_size + 1) downto 0);
        s : out std_logic_vector((total_size - 1) downto 0)
    );
end component;

component adder_compressor_3_2
    Generic(
        total_size : integer
    );
    Port (
        a : in std_logic_vector((total_size - 1) downto 0);
        b : in std_logic_vector((total_size - 1) downto 0);
        p : in std_logic_vector((total_size - 1) downto 0);
        c : out std_logic_vector((total_size) downto 0);
        s : out std_logic_vector((total_size - 1) downto 0)
    );
end component;

component wide_adder_carry_select
    Generic(
        base_size : integer;
        total_size : integer
    );
    Port (
        a : in std_logic_vector((total_size - 1) downto 0);
        b : in std_logic_vector((total_size - 1) downto 0);
        cin : in std_logic_vector(0 downto 0);
        o : out std_logic_vector((total_size - 1) downto 0)
    );
end component;

signal temp_mult_0 : std_logic_vector(40 downto 0);
signal temp_mult_1 : std_logic_vector(64 downto 24);
signal temp_mult_2 : std_logic_vector(88 downto 48);
signal temp_mult_3 : std_logic_vector(112 downto 72);
signal temp_mult_4 : std_logic_vector(136 downto 96);
signal temp_mult_5 : std_logic_vector(57 downto 17);
signal temp_mult_6 : std_logic_vector(81 downto 41);
signal temp_mult_7 : std_logic_vector(105 downto 65);
signal temp_mult_8 : std_logic_vector(129 downto 89);
signal temp_mult_9 : std_logic_vector(153 downto 113);
signal temp_mult_10 : std_logic_vector(74 downto 34);
signal temp_mult_11 : std_logic_vector(98 downto 58);
signal temp_mult_12 : std_logic_vector(122 downto 82);
signal temp_mult_13 : std_logic_vector(146 downto 106);
signal temp_mult_14 : std_logic_vector(170 downto 130);
signal temp_mult_15 : std_logic_vector(91 downto 51);
signal temp_mult_16 : std_logic_vector(115 downto 75);
signal temp_mult_17 : std_logic_vector(139 downto 99);
signal temp_mult_18 : std_logic_vector(163 downto 123);
signal temp_mult_19 : std_logic_vector(187 downto 147);
signal temp_mult_20 : std_logic_vector(108 downto 68);
signal temp_mult_21 : std_logic_vector(132 downto 92);
signal temp_mult_22 : std_logic_vector(156 downto 116);
signal temp_mult_23 : std_logic_vector(180 downto 140);
signal temp_mult_24 : std_logic_vector(204 downto 164);
signal temp_mult_25 : std_logic_vector(125 downto 85);
signal temp_mult_26 : std_logic_vector(149 downto 109);
signal temp_mult_27 : std_logic_vector(173 downto 133);
signal temp_mult_28 : std_logic_vector(197 downto 157);
signal temp_mult_29 : std_logic_vector(221 downto 181);
signal temp_mult_30 : std_logic_vector(142 downto 102);
signal temp_mult_31 : std_logic_vector(166 downto 126);
signal temp_mult_32 : std_logic_vector(190 downto 150);
signal temp_mult_33 : std_logic_vector(214 downto 174);
signal temp_mult_34 : std_logic_vector(238 downto 198);
signal temp_mult_35 : std_logic_vector(159 downto 119);
signal temp_mult_36 : std_logic_vector(183 downto 143);
signal temp_mult_37 : std_logic_vector(207 downto 167);
signal temp_mult_38 : std_logic_vector(231 downto 191);
signal temp_mult_39 : std_logic_vector(255 downto 215);
signal temp_mult_40 : std_logic_vector(160 downto 120);
signal temp_mult_41 : std_logic_vector(177 downto 137);
signal temp_mult_42 : std_logic_vector(194 downto 154);
signal temp_mult_43 : std_logic_vector(211 downto 171);
signal temp_mult_44 : std_logic_vector(228 downto 188);
signal temp_mult_45 : std_logic_vector(245 downto 205);
signal temp_mult_46 : std_logic_vector(262 downto 222);
signal temp_mult_47 : std_logic_vector(279 downto 239);
signal temp_mult_48 : std_logic_vector(184 downto 144);
signal temp_mult_49 : std_logic_vector(201 downto 161);
signal temp_mult_50 : std_logic_vector(218 downto 178);
signal temp_mult_51 : std_logic_vector(235 downto 195);
signal temp_mult_52 : std_logic_vector(252 downto 212);
signal temp_mult_53 : std_logic_vector(269 downto 229);
signal temp_mult_54 : std_logic_vector(286 downto 246);
signal temp_mult_55 : std_logic_vector(303 downto 263);
signal temp_mult_56 : std_logic_vector(208 downto 168);
signal temp_mult_57 : std_logic_vector(225 downto 185);
signal temp_mult_58 : std_logic_vector(242 downto 202);
signal temp_mult_59 : std_logic_vector(259 downto 219);
signal temp_mult_60 : std_logic_vector(276 downto 236);
signal temp_mult_61 : std_logic_vector(293 downto 253);
signal temp_mult_62 : std_logic_vector(310 downto 270);
signal temp_mult_63 : std_logic_vector(327 downto 287);
signal temp_mult_64 : std_logic_vector(232 downto 192);
signal temp_mult_65 : std_logic_vector(249 downto 209);
signal temp_mult_66 : std_logic_vector(266 downto 226);
signal temp_mult_67 : std_logic_vector(283 downto 243);
signal temp_mult_68 : std_logic_vector(300 downto 260);
signal temp_mult_69 : std_logic_vector(317 downto 277);
signal temp_mult_70 : std_logic_vector(334 downto 294);
signal temp_mult_71 : std_logic_vector(351 downto 311);
signal temp_mult_72 : std_logic_vector(256 downto 216);
signal temp_mult_73 : std_logic_vector(273 downto 233);
signal temp_mult_74 : std_logic_vector(290 downto 250);
signal temp_mult_75 : std_logic_vector(307 downto 267);
signal temp_mult_76 : std_logic_vector(324 downto 284);
signal temp_mult_77 : std_logic_vector(341 downto 301);
signal temp_mult_78 : std_logic_vector(358 downto 318);
signal temp_mult_79 : std_logic_vector(375 downto 335);
signal temp_mult_80 : std_logic_vector(176 downto 136);
signal temp_mult_81 : std_logic_vector(193 downto 153);
signal temp_mult_82 : std_logic_vector(210 downto 170);
signal temp_mult_83 : std_logic_vector(227 downto 187);
signal temp_mult_84 : std_logic_vector(244 downto 204);
signal temp_mult_85 : std_logic_vector(261 downto 221);
signal temp_mult_86 : std_logic_vector(278 downto 238);
signal temp_mult_87 : std_logic_vector(295 downto 255);
signal temp_mult_88 : std_logic_vector(200 downto 160);
signal temp_mult_89 : std_logic_vector(217 downto 177);
signal temp_mult_90 : std_logic_vector(234 downto 194);
signal temp_mult_91 : std_logic_vector(251 downto 211);
signal temp_mult_92 : std_logic_vector(268 downto 228);
signal temp_mult_93 : std_logic_vector(285 downto 245);
signal temp_mult_94 : std_logic_vector(302 downto 262);
signal temp_mult_95 : std_logic_vector(319 downto 279);
signal temp_mult_96 : std_logic_vector(224 downto 184);
signal temp_mult_97 : std_logic_vector(241 downto 201);
signal temp_mult_98 : std_logic_vector(258 downto 218);
signal temp_mult_99 : std_logic_vector(275 downto 235);
signal temp_mult_100 : std_logic_vector(292 downto 252);
signal temp_mult_101 : std_logic_vector(309 downto 269);
signal temp_mult_102 : std_logic_vector(326 downto 286);
signal temp_mult_103 : std_logic_vector(343 downto 303);
signal temp_mult_104 : std_logic_vector(248 downto 208);
signal temp_mult_105 : std_logic_vector(265 downto 225);
signal temp_mult_106 : std_logic_vector(282 downto 242);
signal temp_mult_107 : std_logic_vector(299 downto 259);
signal temp_mult_108 : std_logic_vector(316 downto 276);
signal temp_mult_109 : std_logic_vector(333 downto 293);
signal temp_mult_110 : std_logic_vector(350 downto 310);
signal temp_mult_111 : std_logic_vector(367 downto 327);
signal temp_mult_112 : std_logic_vector(272 downto 232);
signal temp_mult_113 : std_logic_vector(289 downto 249);
signal temp_mult_114 : std_logic_vector(306 downto 266);
signal temp_mult_115 : std_logic_vector(323 downto 283);
signal temp_mult_116 : std_logic_vector(340 downto 300);
signal temp_mult_117 : std_logic_vector(357 downto 317);
signal temp_mult_118 : std_logic_vector(374 downto 334);
signal temp_mult_119 : std_logic_vector(391 downto 351);
signal temp_mult_120 : std_logic_vector(296 downto 256);
signal temp_mult_121 : std_logic_vector(320 downto 280);
signal temp_mult_122 : std_logic_vector(344 downto 304);
signal temp_mult_123 : std_logic_vector(368 downto 328);
signal temp_mult_124 : std_logic_vector(392 downto 352);
signal temp_mult_125 : std_logic_vector(313 downto 273);
signal temp_mult_126 : std_logic_vector(337 downto 297);
signal temp_mult_127 : std_logic_vector(361 downto 321);
signal temp_mult_128 : std_logic_vector(385 downto 345);
signal temp_mult_129 : std_logic_vector(409 downto 369);
signal temp_mult_130 : std_logic_vector(330 downto 290);
signal temp_mult_131 : std_logic_vector(354 downto 314);
signal temp_mult_132 : std_logic_vector(378 downto 338);
signal temp_mult_133 : std_logic_vector(402 downto 362);
signal temp_mult_134 : std_logic_vector(426 downto 386);
signal temp_mult_135 : std_logic_vector(347 downto 307);
signal temp_mult_136 : std_logic_vector(371 downto 331);
signal temp_mult_137 : std_logic_vector(395 downto 355);
signal temp_mult_138 : std_logic_vector(419 downto 379);
signal temp_mult_139 : std_logic_vector(443 downto 403);
signal temp_mult_140 : std_logic_vector(364 downto 324);
signal temp_mult_141 : std_logic_vector(388 downto 348);
signal temp_mult_142 : std_logic_vector(412 downto 372);
signal temp_mult_143 : std_logic_vector(436 downto 396);
signal temp_mult_144 : std_logic_vector(460 downto 420);
signal temp_mult_145 : std_logic_vector(381 downto 341);
signal temp_mult_146 : std_logic_vector(405 downto 365);
signal temp_mult_147 : std_logic_vector(429 downto 389);
signal temp_mult_148 : std_logic_vector(453 downto 413);
signal temp_mult_149 : std_logic_vector(477 downto 437);
signal temp_mult_150 : std_logic_vector(398 downto 358);
signal temp_mult_151 : std_logic_vector(422 downto 382);
signal temp_mult_152 : std_logic_vector(446 downto 406);
signal temp_mult_153 : std_logic_vector(470 downto 430);
signal temp_mult_154 : std_logic_vector(494 downto 454);
signal temp_mult_155 : std_logic_vector(415 downto 375);
signal temp_mult_156 : std_logic_vector(439 downto 399);
signal temp_mult_157 : std_logic_vector(463 downto 423);
signal temp_mult_158 : std_logic_vector(487 downto 447);
signal temp_mult_159 : std_logic_vector(511 downto 471);
signal temp_mult_160 : std_logic_vector(271 downto 240);
signal temp_part_mult_161 : std_logic_vector(511 downto 256);
signal temp_part_mult_162 : std_logic_vector(512 downto 256);
signal temp_mult_161 : std_logic_vector(513 downto 256);
signal temp_mult_162 : std_logic_vector(513 downto 256);

signal partial_product_0 : std_logic_vector(512 downto 0);
signal partial_product_1 : std_logic_vector(512 downto 0);
signal partial_product_2 : std_logic_vector(512 downto 0);
signal partial_product_3 : std_logic_vector(512 downto 0);
signal partial_product_4 : std_logic_vector(512 downto 0);
signal partial_product_5 : std_logic_vector(512 downto 0);
signal partial_product_6 : std_logic_vector(512 downto 0);
signal partial_product_7 : std_logic_vector(512 downto 0);
signal partial_product_8 : std_logic_vector(512 downto 0);
signal partial_product_9 : std_logic_vector(512 downto 0);
signal partial_product_10 : std_logic_vector(512 downto 0);
signal partial_product_11 : std_logic_vector(512 downto 0);
signal partial_product_12 : std_logic_vector(512 downto 0);
signal partial_product_13 : std_logic_vector(512 downto 0);
signal partial_product_14 : std_logic_vector(512 downto 0);
signal partial_product_15 : std_logic_vector(512 downto 0);
signal partial_product_16 : std_logic_vector(512 downto 0);
signal partial_product_17 : std_logic_vector(512 downto 0);
signal partial_product_18 : std_logic_vector(512 downto 0);
signal partial_product_19 : std_logic_vector(512 downto 0);
signal partial_product_20 : std_logic_vector(512 downto 0);
signal partial_product_21 : std_logic_vector(512 downto 0);
signal partial_product_22 : std_logic_vector(512 downto 0);
signal partial_product_23 : std_logic_vector(512 downto 0);
signal partial_product_24 : std_logic_vector(512 downto 0);
signal partial_product_25 : std_logic_vector(512 downto 0);
signal partial_product_26 : std_logic_vector(513 downto 0);
signal partial_product_27 : std_logic_vector(513 downto 0);

signal temp_comp_1_a1 : std_logic_vector(513 downto 0);
signal temp_comp_1_a2 : std_logic_vector(513 downto 0);
signal temp_comp_1_a3 : std_logic_vector(513 downto 0);
signal temp_comp_1_a4 : std_logic_vector(513 downto 0);
signal temp_comp_1_a5 : std_logic_vector(513 downto 0);
signal temp_comp_1_a6 : std_logic_vector(513 downto 0);
signal temp_comp_1_a7 : std_logic_vector(513 downto 0);
signal temp_comp_1_a8 : std_logic_vector(513 downto 0);
signal temp_comp_1_a9 : std_logic_vector(513 downto 0);
signal temp_comp_1_a10 : std_logic_vector(513 downto 0);
signal temp_comp_1_a11 : std_logic_vector(513 downto 0);
signal temp_comp_1_a12 : std_logic_vector(513 downto 0);
signal temp_comp_1_a13 : std_logic_vector(513 downto 0);
signal temp_comp_1_a14 : std_logic_vector(513 downto 0);
signal temp_comp_1_a15 : std_logic_vector(513 downto 0);
signal temp_comp_1_a16 : std_logic_vector(513 downto 0);
signal temp_comp_1_a17 : std_logic_vector(513 downto 0);
signal temp_comp_1_a18 : std_logic_vector(513 downto 0);
signal temp_comp_1_a19 : std_logic_vector(513 downto 0);
signal temp_comp_1_a20 : std_logic_vector(513 downto 0);
signal temp_comp_1_a21 : std_logic_vector(513 downto 0);
signal temp_comp_1_a22 : std_logic_vector(513 downto 0);
signal temp_comp_1_a23 : std_logic_vector(513 downto 0);
signal temp_comp_1_a24 : std_logic_vector(513 downto 0);
signal temp_comp_1_a25 : std_logic_vector(513 downto 0);
signal temp_comp_1_a26 : std_logic_vector(513 downto 0);
signal temp_comp_1_a27 : std_logic_vector(513 downto 0);
signal temp_comp_1_a28 : std_logic_vector(513 downto 0);
signal temp_comp_1_a29 : std_logic_vector(513 downto 0);
signal temp_comp_1_a30 : std_logic_vector(513 downto 0);
signal temp_comp_1_c1 : std_logic_vector(514 downto 0);
signal temp_comp_1_c2 : std_logic_vector(515 downto 0);
signal temp_comp_1_c3 : std_logic_vector(516 downto 0);
signal temp_comp_1_c4 : std_logic_vector(517 downto 0);
signal temp_comp_1_s : std_logic_vector(513 downto 0);

signal temp_comp_2_a1 : std_logic_vector(513 downto 0);
signal temp_comp_2_a2 : std_logic_vector(513 downto 0);
signal temp_comp_2_a3 : std_logic_vector(513 downto 0);
signal temp_comp_2_a4 : std_logic_vector(513 downto 0);
signal temp_comp_2_a5 : std_logic_vector(513 downto 0);
signal temp_comp_2_c1 : std_logic_vector(514 downto 0);
signal temp_comp_2_c2 : std_logic_vector(515 downto 0);
signal temp_comp_2_s : std_logic_vector(513 downto 0);

signal temp_comp_3_a1 : std_logic_vector(513 downto 0);
signal temp_comp_3_a2 : std_logic_vector(513 downto 0);
signal temp_comp_3_a3 : std_logic_vector(513 downto 0);
signal temp_comp_3_c  : std_logic_vector(514 downto 0);
signal temp_comp_3_s  : std_logic_vector(513 downto 0);

signal temp_comp_4_a1 : std_logic_vector(513 downto 0);
signal temp_comp_4_a2 : std_logic_vector(513 downto 0);

signal final_comp_a : std_logic_vector(513 downto 0);
signal final_comp_b : std_logic_vector(513 downto 0);
signal final_comp_o : std_logic_vector(513 downto 0);

signal temp_o4 : unsigned(513 downto 0);
signal temp_o5 : unsigned(513 downto 0);


begin

temp_mult_0 <= std_logic_vector(unsigned(a(16 downto 0)) * unsigned(b(23 downto 0))); 
temp_mult_1 <= std_logic_vector(unsigned(a(16 downto 0)) * unsigned(b(47 downto 24))); 
temp_mult_2 <= std_logic_vector(unsigned(a(16 downto 0)) * unsigned(b(71 downto 48))); 
temp_mult_3 <= std_logic_vector(unsigned(a(16 downto 0)) * unsigned(b(95 downto 72))); 
temp_mult_4 <= std_logic_vector(unsigned(a(16 downto 0)) * unsigned(b(119 downto 96))); 
temp_mult_5 <= std_logic_vector(unsigned(a(33 downto 17)) * unsigned(b(23 downto 0))); 
temp_mult_6 <= std_logic_vector(unsigned(a(33 downto 17)) * unsigned(b(47 downto 24))); 
temp_mult_7 <= std_logic_vector(unsigned(a(33 downto 17)) * unsigned(b(71 downto 48))); 
temp_mult_8 <= std_logic_vector(unsigned(a(33 downto 17)) * unsigned(b(95 downto 72))); 
temp_mult_9 <= std_logic_vector(unsigned(a(33 downto 17)) * unsigned(b(119 downto 96))); 
temp_mult_10 <= std_logic_vector(unsigned(a(50 downto 34)) * unsigned(b(23 downto 0))); 
temp_mult_11 <= std_logic_vector(unsigned(a(50 downto 34)) * unsigned(b(47 downto 24))); 
temp_mult_12 <= std_logic_vector(unsigned(a(50 downto 34)) * unsigned(b(71 downto 48))); 
temp_mult_13 <= std_logic_vector(unsigned(a(50 downto 34)) * unsigned(b(95 downto 72))); 
temp_mult_14 <= std_logic_vector(unsigned(a(50 downto 34)) * unsigned(b(119 downto 96))); 
temp_mult_15 <= std_logic_vector(unsigned(a(67 downto 51)) * unsigned(b(23 downto 0))); 
temp_mult_16 <= std_logic_vector(unsigned(a(67 downto 51)) * unsigned(b(47 downto 24))); 
temp_mult_17 <= std_logic_vector(unsigned(a(67 downto 51)) * unsigned(b(71 downto 48))); 
temp_mult_18 <= std_logic_vector(unsigned(a(67 downto 51)) * unsigned(b(95 downto 72))); 
temp_mult_19 <= std_logic_vector(unsigned(a(67 downto 51)) * unsigned(b(119 downto 96))); 
temp_mult_20 <= std_logic_vector(unsigned(a(84 downto 68)) * unsigned(b(23 downto 0))); 
temp_mult_21 <= std_logic_vector(unsigned(a(84 downto 68)) * unsigned(b(47 downto 24))); 
temp_mult_22 <= std_logic_vector(unsigned(a(84 downto 68)) * unsigned(b(71 downto 48))); 
temp_mult_23 <= std_logic_vector(unsigned(a(84 downto 68)) * unsigned(b(95 downto 72))); 
temp_mult_24 <= std_logic_vector(unsigned(a(84 downto 68)) * unsigned(b(119 downto 96))); 
temp_mult_25 <= std_logic_vector(unsigned(a(101 downto 85)) * unsigned(b(23 downto 0))); 
temp_mult_26 <= std_logic_vector(unsigned(a(101 downto 85)) * unsigned(b(47 downto 24))); 
temp_mult_27 <= std_logic_vector(unsigned(a(101 downto 85)) * unsigned(b(71 downto 48))); 
temp_mult_28 <= std_logic_vector(unsigned(a(101 downto 85)) * unsigned(b(95 downto 72))); 
temp_mult_29 <= std_logic_vector(unsigned(a(101 downto 85)) * unsigned(b(119 downto 96))); 
temp_mult_30 <= std_logic_vector(unsigned(a(118 downto 102)) * unsigned(b(23 downto 0))); 
temp_mult_31 <= std_logic_vector(unsigned(a(118 downto 102)) * unsigned(b(47 downto 24))); 
temp_mult_32 <= std_logic_vector(unsigned(a(118 downto 102)) * unsigned(b(71 downto 48))); 
temp_mult_33 <= std_logic_vector(unsigned(a(118 downto 102)) * unsigned(b(95 downto 72))); 
temp_mult_34 <= std_logic_vector(unsigned(a(118 downto 102)) * unsigned(b(119 downto 96))); 
temp_mult_35 <= std_logic_vector(unsigned(a(135 downto 119)) * unsigned(b(23 downto 0))); 
temp_mult_36 <= std_logic_vector(unsigned(a(135 downto 119)) * unsigned(b(47 downto 24))); 
temp_mult_37 <= std_logic_vector(unsigned(a(135 downto 119)) * unsigned(b(71 downto 48))); 
temp_mult_38 <= std_logic_vector(unsigned(a(135 downto 119)) * unsigned(b(95 downto 72))); 
temp_mult_39 <= std_logic_vector(unsigned(a(135 downto 119)) * unsigned(b(119 downto 96))); 
temp_mult_40 <= std_logic_vector(unsigned(a(23 downto 0)) * unsigned(b(136 downto 120))); 
temp_mult_41 <= std_logic_vector(unsigned(a(23 downto 0)) * unsigned(b(153 downto 137))); 
temp_mult_42 <= std_logic_vector(unsigned(a(23 downto 0)) * unsigned(b(170 downto 154))); 
temp_mult_43 <= std_logic_vector(unsigned(a(23 downto 0)) * unsigned(b(187 downto 171))); 
temp_mult_44 <= std_logic_vector(unsigned(a(23 downto 0)) * unsigned(b(204 downto 188))); 
temp_mult_45 <= std_logic_vector(unsigned(a(23 downto 0)) * unsigned(b(221 downto 205))); 
temp_mult_46 <= std_logic_vector(unsigned(a(23 downto 0)) * unsigned(b(238 downto 222))); 
temp_mult_47 <= std_logic_vector(unsigned(a(23 downto 0)) * unsigned(b(255 downto 239))); 
temp_mult_48 <= std_logic_vector(unsigned(a(47 downto 24)) * unsigned(b(136 downto 120))); 
temp_mult_49 <= std_logic_vector(unsigned(a(47 downto 24)) * unsigned(b(153 downto 137))); 
temp_mult_50 <= std_logic_vector(unsigned(a(47 downto 24)) * unsigned(b(170 downto 154))); 
temp_mult_51 <= std_logic_vector(unsigned(a(47 downto 24)) * unsigned(b(187 downto 171))); 
temp_mult_52 <= std_logic_vector(unsigned(a(47 downto 24)) * unsigned(b(204 downto 188))); 
temp_mult_53 <= std_logic_vector(unsigned(a(47 downto 24)) * unsigned(b(221 downto 205))); 
temp_mult_54 <= std_logic_vector(unsigned(a(47 downto 24)) * unsigned(b(238 downto 222))); 
temp_mult_55 <= std_logic_vector(unsigned(a(47 downto 24)) * unsigned(b(255 downto 239))); 
temp_mult_56 <= std_logic_vector(unsigned(a(71 downto 48)) * unsigned(b(136 downto 120))); 
temp_mult_57 <= std_logic_vector(unsigned(a(71 downto 48)) * unsigned(b(153 downto 137))); 
temp_mult_58 <= std_logic_vector(unsigned(a(71 downto 48)) * unsigned(b(170 downto 154))); 
temp_mult_59 <= std_logic_vector(unsigned(a(71 downto 48)) * unsigned(b(187 downto 171))); 
temp_mult_60 <= std_logic_vector(unsigned(a(71 downto 48)) * unsigned(b(204 downto 188))); 
temp_mult_61 <= std_logic_vector(unsigned(a(71 downto 48)) * unsigned(b(221 downto 205))); 
temp_mult_62 <= std_logic_vector(unsigned(a(71 downto 48)) * unsigned(b(238 downto 222))); 
temp_mult_63 <= std_logic_vector(unsigned(a(71 downto 48)) * unsigned(b(255 downto 239))); 
temp_mult_64 <= std_logic_vector(unsigned(a(95 downto 72)) * unsigned(b(136 downto 120))); 
temp_mult_65 <= std_logic_vector(unsigned(a(95 downto 72)) * unsigned(b(153 downto 137))); 
temp_mult_66 <= std_logic_vector(unsigned(a(95 downto 72)) * unsigned(b(170 downto 154))); 
temp_mult_67 <= std_logic_vector(unsigned(a(95 downto 72)) * unsigned(b(187 downto 171))); 
temp_mult_68 <= std_logic_vector(unsigned(a(95 downto 72)) * unsigned(b(204 downto 188))); 
temp_mult_69 <= std_logic_vector(unsigned(a(95 downto 72)) * unsigned(b(221 downto 205))); 
temp_mult_70 <= std_logic_vector(unsigned(a(95 downto 72)) * unsigned(b(238 downto 222))); 
temp_mult_71 <= std_logic_vector(unsigned(a(95 downto 72)) * unsigned(b(255 downto 239))); 
temp_mult_72 <= std_logic_vector(unsigned(a(119 downto 96)) * unsigned(b(136 downto 120))); 
temp_mult_73 <= std_logic_vector(unsigned(a(119 downto 96)) * unsigned(b(153 downto 137))); 
temp_mult_74 <= std_logic_vector(unsigned(a(119 downto 96)) * unsigned(b(170 downto 154))); 
temp_mult_75 <= std_logic_vector(unsigned(a(119 downto 96)) * unsigned(b(187 downto 171))); 
temp_mult_76 <= std_logic_vector(unsigned(a(119 downto 96)) * unsigned(b(204 downto 188))); 
temp_mult_77 <= std_logic_vector(unsigned(a(119 downto 96)) * unsigned(b(221 downto 205))); 
temp_mult_78 <= std_logic_vector(unsigned(a(119 downto 96)) * unsigned(b(238 downto 222))); 
temp_mult_79 <= std_logic_vector(unsigned(a(119 downto 96)) * unsigned(b(255 downto 239))); 
temp_mult_80 <= std_logic_vector(unsigned(a(159 downto 136)) * unsigned(b(16 downto 0))); 
temp_mult_81 <= std_logic_vector(unsigned(a(159 downto 136)) * unsigned(b(33 downto 17))); 
temp_mult_82 <= std_logic_vector(unsigned(a(159 downto 136)) * unsigned(b(50 downto 34))); 
temp_mult_83 <= std_logic_vector(unsigned(a(159 downto 136)) * unsigned(b(67 downto 51))); 
temp_mult_84 <= std_logic_vector(unsigned(a(159 downto 136)) * unsigned(b(84 downto 68))); 
temp_mult_85 <= std_logic_vector(unsigned(a(159 downto 136)) * unsigned(b(101 downto 85))); 
temp_mult_86 <= std_logic_vector(unsigned(a(159 downto 136)) * unsigned(b(118 downto 102))); 
temp_mult_87 <= std_logic_vector(unsigned(a(159 downto 136)) * unsigned(b(135 downto 119))); 
temp_mult_88 <= std_logic_vector(unsigned(a(183 downto 160)) * unsigned(b(16 downto 0))); 
temp_mult_89 <= std_logic_vector(unsigned(a(183 downto 160)) * unsigned(b(33 downto 17))); 
temp_mult_90 <= std_logic_vector(unsigned(a(183 downto 160)) * unsigned(b(50 downto 34))); 
temp_mult_91 <= std_logic_vector(unsigned(a(183 downto 160)) * unsigned(b(67 downto 51))); 
temp_mult_92 <= std_logic_vector(unsigned(a(183 downto 160)) * unsigned(b(84 downto 68))); 
temp_mult_93 <= std_logic_vector(unsigned(a(183 downto 160)) * unsigned(b(101 downto 85))); 
temp_mult_94 <= std_logic_vector(unsigned(a(183 downto 160)) * unsigned(b(118 downto 102))); 
temp_mult_95 <= std_logic_vector(unsigned(a(183 downto 160)) * unsigned(b(135 downto 119))); 
temp_mult_96 <= std_logic_vector(unsigned(a(207 downto 184)) * unsigned(b(16 downto 0))); 
temp_mult_97 <= std_logic_vector(unsigned(a(207 downto 184)) * unsigned(b(33 downto 17))); 
temp_mult_98 <= std_logic_vector(unsigned(a(207 downto 184)) * unsigned(b(50 downto 34))); 
temp_mult_99 <= std_logic_vector(unsigned(a(207 downto 184)) * unsigned(b(67 downto 51))); 
temp_mult_100 <= std_logic_vector(unsigned(a(207 downto 184)) * unsigned(b(84 downto 68))); 
temp_mult_101 <= std_logic_vector(unsigned(a(207 downto 184)) * unsigned(b(101 downto 85))); 
temp_mult_102 <= std_logic_vector(unsigned(a(207 downto 184)) * unsigned(b(118 downto 102))); 
temp_mult_103 <= std_logic_vector(unsigned(a(207 downto 184)) * unsigned(b(135 downto 119))); 
temp_mult_104 <= std_logic_vector(unsigned(a(231 downto 208)) * unsigned(b(16 downto 0))); 
temp_mult_105 <= std_logic_vector(unsigned(a(231 downto 208)) * unsigned(b(33 downto 17))); 
temp_mult_106 <= std_logic_vector(unsigned(a(231 downto 208)) * unsigned(b(50 downto 34))); 
temp_mult_107 <= std_logic_vector(unsigned(a(231 downto 208)) * unsigned(b(67 downto 51))); 
temp_mult_108 <= std_logic_vector(unsigned(a(231 downto 208)) * unsigned(b(84 downto 68))); 
temp_mult_109 <= std_logic_vector(unsigned(a(231 downto 208)) * unsigned(b(101 downto 85))); 
temp_mult_110 <= std_logic_vector(unsigned(a(231 downto 208)) * unsigned(b(118 downto 102))); 
temp_mult_111 <= std_logic_vector(unsigned(a(231 downto 208)) * unsigned(b(135 downto 119))); 
temp_mult_112 <= std_logic_vector(unsigned(a(255 downto 232)) * unsigned(b(16 downto 0))); 
temp_mult_113 <= std_logic_vector(unsigned(a(255 downto 232)) * unsigned(b(33 downto 17))); 
temp_mult_114 <= std_logic_vector(unsigned(a(255 downto 232)) * unsigned(b(50 downto 34))); 
temp_mult_115 <= std_logic_vector(unsigned(a(255 downto 232)) * unsigned(b(67 downto 51))); 
temp_mult_116 <= std_logic_vector(unsigned(a(255 downto 232)) * unsigned(b(84 downto 68))); 
temp_mult_117 <= std_logic_vector(unsigned(a(255 downto 232)) * unsigned(b(101 downto 85))); 
temp_mult_118 <= std_logic_vector(unsigned(a(255 downto 232)) * unsigned(b(118 downto 102))); 
temp_mult_119 <= std_logic_vector(unsigned(a(255 downto 232)) * unsigned(b(135 downto 119))); 
temp_mult_120 <= std_logic_vector(unsigned(a(136 downto 120)) * unsigned(b(159 downto 136))); 
temp_mult_121 <= std_logic_vector(unsigned(a(136 downto 120)) * unsigned(b(183 downto 160))); 
temp_mult_122 <= std_logic_vector(unsigned(a(136 downto 120)) * unsigned(b(207 downto 184))); 
temp_mult_123 <= std_logic_vector(unsigned(a(136 downto 120)) * unsigned(b(231 downto 208))); 
temp_mult_124 <= std_logic_vector(unsigned(a(136 downto 120)) * unsigned(b(255 downto 232))); 
temp_mult_125 <= std_logic_vector(unsigned(a(153 downto 137)) * unsigned(b(159 downto 136))); 
temp_mult_126 <= std_logic_vector(unsigned(a(153 downto 137)) * unsigned(b(183 downto 160))); 
temp_mult_127 <= std_logic_vector(unsigned(a(153 downto 137)) * unsigned(b(207 downto 184))); 
temp_mult_128 <= std_logic_vector(unsigned(a(153 downto 137)) * unsigned(b(231 downto 208))); 
temp_mult_129 <= std_logic_vector(unsigned(a(153 downto 137)) * unsigned(b(255 downto 232))); 
temp_mult_130 <= std_logic_vector(unsigned(a(170 downto 154)) * unsigned(b(159 downto 136))); 
temp_mult_131 <= std_logic_vector(unsigned(a(170 downto 154)) * unsigned(b(183 downto 160))); 
temp_mult_132 <= std_logic_vector(unsigned(a(170 downto 154)) * unsigned(b(207 downto 184))); 
temp_mult_133 <= std_logic_vector(unsigned(a(170 downto 154)) * unsigned(b(231 downto 208))); 
temp_mult_134 <= std_logic_vector(unsigned(a(170 downto 154)) * unsigned(b(255 downto 232))); 
temp_mult_135 <= std_logic_vector(unsigned(a(187 downto 171)) * unsigned(b(159 downto 136))); 
temp_mult_136 <= std_logic_vector(unsigned(a(187 downto 171)) * unsigned(b(183 downto 160))); 
temp_mult_137 <= std_logic_vector(unsigned(a(187 downto 171)) * unsigned(b(207 downto 184))); 
temp_mult_138 <= std_logic_vector(unsigned(a(187 downto 171)) * unsigned(b(231 downto 208))); 
temp_mult_139 <= std_logic_vector(unsigned(a(187 downto 171)) * unsigned(b(255 downto 232))); 
temp_mult_140 <= std_logic_vector(unsigned(a(204 downto 188)) * unsigned(b(159 downto 136))); 
temp_mult_141 <= std_logic_vector(unsigned(a(204 downto 188)) * unsigned(b(183 downto 160))); 
temp_mult_142 <= std_logic_vector(unsigned(a(204 downto 188)) * unsigned(b(207 downto 184))); 
temp_mult_143 <= std_logic_vector(unsigned(a(204 downto 188)) * unsigned(b(231 downto 208))); 
temp_mult_144 <= std_logic_vector(unsigned(a(204 downto 188)) * unsigned(b(255 downto 232))); 
temp_mult_145 <= std_logic_vector(unsigned(a(221 downto 205)) * unsigned(b(159 downto 136))); 
temp_mult_146 <= std_logic_vector(unsigned(a(221 downto 205)) * unsigned(b(183 downto 160))); 
temp_mult_147 <= std_logic_vector(unsigned(a(221 downto 205)) * unsigned(b(207 downto 184))); 
temp_mult_148 <= std_logic_vector(unsigned(a(221 downto 205)) * unsigned(b(231 downto 208))); 
temp_mult_149 <= std_logic_vector(unsigned(a(221 downto 205)) * unsigned(b(255 downto 232))); 
temp_mult_150 <= std_logic_vector(unsigned(a(238 downto 222)) * unsigned(b(159 downto 136))); 
temp_mult_151 <= std_logic_vector(unsigned(a(238 downto 222)) * unsigned(b(183 downto 160))); 
temp_mult_152 <= std_logic_vector(unsigned(a(238 downto 222)) * unsigned(b(207 downto 184))); 
temp_mult_153 <= std_logic_vector(unsigned(a(238 downto 222)) * unsigned(b(231 downto 208))); 
temp_mult_154 <= std_logic_vector(unsigned(a(238 downto 222)) * unsigned(b(255 downto 232))); 
temp_mult_155 <= std_logic_vector(unsigned(a(255 downto 239)) * unsigned(b(159 downto 136))); 
temp_mult_156 <= std_logic_vector(unsigned(a(255 downto 239)) * unsigned(b(183 downto 160))); 
temp_mult_157 <= std_logic_vector(unsigned(a(255 downto 239)) * unsigned(b(207 downto 184))); 
temp_mult_158 <= std_logic_vector(unsigned(a(255 downto 239)) * unsigned(b(231 downto 208))); 
temp_mult_159 <= std_logic_vector(unsigned(a(255 downto 239)) * unsigned(b(255 downto 232))); 
temp_mult_160 <= std_logic_vector(unsigned(a(135 downto 120)) * unsigned(b(135 downto 120))); 
temp_part_mult_161 <= (others => a(256));
temp_part_mult_162 <= (others => b(256));
temp_mult_161(511 downto 256) <= temp_part_mult_161 and b(255 downto 0);
temp_mult_161(513 downto 512) <= "00";
temp_mult_162(512 downto 256) <= temp_part_mult_162 and a(256 downto 0); 
temp_mult_162(513) <= temp_mult_162(512); 

partial_product_0(0) <= temp_mult_0(0);
partial_product_0(1) <= temp_mult_0(1);
partial_product_0(2) <= temp_mult_0(2);
partial_product_0(3) <= temp_mult_0(3);
partial_product_0(4) <= temp_mult_0(4);
partial_product_0(5) <= temp_mult_0(5);
partial_product_0(6) <= temp_mult_0(6);
partial_product_0(7) <= temp_mult_0(7);
partial_product_0(8) <= temp_mult_0(8);
partial_product_0(9) <= temp_mult_0(9);
partial_product_0(10) <= temp_mult_0(10);
partial_product_0(11) <= temp_mult_0(11);
partial_product_0(12) <= temp_mult_0(12);
partial_product_0(13) <= temp_mult_0(13);
partial_product_0(14) <= temp_mult_0(14);
partial_product_0(15) <= temp_mult_0(15);
partial_product_0(16) <= temp_mult_0(16);
partial_product_0(17) <= temp_mult_0(17);
partial_product_0(18) <= temp_mult_0(18);
partial_product_0(19) <= temp_mult_0(19);
partial_product_0(20) <= temp_mult_0(20);
partial_product_0(21) <= temp_mult_0(21);
partial_product_0(22) <= temp_mult_0(22);
partial_product_0(23) <= temp_mult_0(23);
partial_product_0(24) <= temp_mult_0(24);
partial_product_0(25) <= temp_mult_0(25);
partial_product_0(26) <= temp_mult_0(26);
partial_product_0(27) <= temp_mult_0(27);
partial_product_0(28) <= temp_mult_0(28);
partial_product_0(29) <= temp_mult_0(29);
partial_product_0(30) <= temp_mult_0(30);
partial_product_0(31) <= temp_mult_0(31);
partial_product_0(32) <= temp_mult_0(32);
partial_product_0(33) <= temp_mult_0(33);
partial_product_0(34) <= temp_mult_0(34);
partial_product_0(35) <= temp_mult_0(35);
partial_product_0(36) <= temp_mult_0(36);
partial_product_0(37) <= temp_mult_0(37);
partial_product_0(38) <= temp_mult_0(38);
partial_product_0(39) <= temp_mult_0(39);
partial_product_0(40) <= temp_mult_0(40);
partial_product_0(41) <= temp_mult_6(41);
partial_product_0(42) <= temp_mult_6(42);
partial_product_0(43) <= temp_mult_6(43);
partial_product_0(44) <= temp_mult_6(44);
partial_product_0(45) <= temp_mult_6(45);
partial_product_0(46) <= temp_mult_6(46);
partial_product_0(47) <= temp_mult_6(47);
partial_product_0(48) <= temp_mult_6(48);
partial_product_0(49) <= temp_mult_6(49);
partial_product_0(50) <= temp_mult_6(50);
partial_product_0(51) <= temp_mult_6(51);
partial_product_0(52) <= temp_mult_6(52);
partial_product_0(53) <= temp_mult_6(53);
partial_product_0(54) <= temp_mult_6(54);
partial_product_0(55) <= temp_mult_6(55);
partial_product_0(56) <= temp_mult_6(56);
partial_product_0(57) <= temp_mult_6(57);
partial_product_0(58) <= temp_mult_6(58);
partial_product_0(59) <= temp_mult_6(59);
partial_product_0(60) <= temp_mult_6(60);
partial_product_0(61) <= temp_mult_6(61);
partial_product_0(62) <= temp_mult_6(62);
partial_product_0(63) <= temp_mult_6(63);
partial_product_0(64) <= temp_mult_6(64);
partial_product_0(65) <= temp_mult_6(65);
partial_product_0(66) <= temp_mult_6(66);
partial_product_0(67) <= temp_mult_6(67);
partial_product_0(68) <= temp_mult_6(68);
partial_product_0(69) <= temp_mult_6(69);
partial_product_0(70) <= temp_mult_6(70);
partial_product_0(71) <= temp_mult_6(71);
partial_product_0(72) <= temp_mult_6(72);
partial_product_0(73) <= temp_mult_6(73);
partial_product_0(74) <= temp_mult_6(74);
partial_product_0(75) <= temp_mult_6(75);
partial_product_0(76) <= temp_mult_6(76);
partial_product_0(77) <= temp_mult_6(77);
partial_product_0(78) <= temp_mult_6(78);
partial_product_0(79) <= temp_mult_6(79);
partial_product_0(80) <= temp_mult_6(80);
partial_product_0(81) <= temp_mult_6(81);
partial_product_0(82) <= temp_mult_12(82);
partial_product_0(83) <= temp_mult_12(83);
partial_product_0(84) <= temp_mult_12(84);
partial_product_0(85) <= temp_mult_12(85);
partial_product_0(86) <= temp_mult_12(86);
partial_product_0(87) <= temp_mult_12(87);
partial_product_0(88) <= temp_mult_12(88);
partial_product_0(89) <= temp_mult_12(89);
partial_product_0(90) <= temp_mult_12(90);
partial_product_0(91) <= temp_mult_12(91);
partial_product_0(92) <= temp_mult_12(92);
partial_product_0(93) <= temp_mult_12(93);
partial_product_0(94) <= temp_mult_12(94);
partial_product_0(95) <= temp_mult_12(95);
partial_product_0(96) <= temp_mult_12(96);
partial_product_0(97) <= temp_mult_12(97);
partial_product_0(98) <= temp_mult_12(98);
partial_product_0(99) <= temp_mult_12(99);
partial_product_0(100) <= temp_mult_12(100);
partial_product_0(101) <= temp_mult_12(101);
partial_product_0(102) <= temp_mult_12(102);
partial_product_0(103) <= temp_mult_12(103);
partial_product_0(104) <= temp_mult_12(104);
partial_product_0(105) <= temp_mult_12(105);
partial_product_0(106) <= temp_mult_12(106);
partial_product_0(107) <= temp_mult_12(107);
partial_product_0(108) <= temp_mult_12(108);
partial_product_0(109) <= temp_mult_12(109);
partial_product_0(110) <= temp_mult_12(110);
partial_product_0(111) <= temp_mult_12(111);
partial_product_0(112) <= temp_mult_12(112);
partial_product_0(113) <= temp_mult_12(113);
partial_product_0(114) <= temp_mult_12(114);
partial_product_0(115) <= temp_mult_12(115);
partial_product_0(116) <= temp_mult_12(116);
partial_product_0(117) <= temp_mult_12(117);
partial_product_0(118) <= temp_mult_12(118);
partial_product_0(119) <= temp_mult_12(119);
partial_product_0(120) <= temp_mult_12(120);
partial_product_0(121) <= temp_mult_12(121);
partial_product_0(122) <= temp_mult_12(122);
partial_product_0(123) <= temp_mult_18(123);
partial_product_0(124) <= temp_mult_18(124);
partial_product_0(125) <= temp_mult_18(125);
partial_product_0(126) <= temp_mult_18(126);
partial_product_0(127) <= temp_mult_18(127);
partial_product_0(128) <= temp_mult_18(128);
partial_product_0(129) <= temp_mult_18(129);
partial_product_0(130) <= temp_mult_18(130);
partial_product_0(131) <= temp_mult_18(131);
partial_product_0(132) <= temp_mult_18(132);
partial_product_0(133) <= temp_mult_18(133);
partial_product_0(134) <= temp_mult_18(134);
partial_product_0(135) <= temp_mult_18(135);
partial_product_0(136) <= temp_mult_18(136);
partial_product_0(137) <= temp_mult_18(137);
partial_product_0(138) <= temp_mult_18(138);
partial_product_0(139) <= temp_mult_18(139);
partial_product_0(140) <= temp_mult_18(140);
partial_product_0(141) <= temp_mult_18(141);
partial_product_0(142) <= temp_mult_18(142);
partial_product_0(143) <= temp_mult_18(143);
partial_product_0(144) <= temp_mult_18(144);
partial_product_0(145) <= temp_mult_18(145);
partial_product_0(146) <= temp_mult_18(146);
partial_product_0(147) <= temp_mult_18(147);
partial_product_0(148) <= temp_mult_18(148);
partial_product_0(149) <= temp_mult_18(149);
partial_product_0(150) <= temp_mult_18(150);
partial_product_0(151) <= temp_mult_18(151);
partial_product_0(152) <= temp_mult_18(152);
partial_product_0(153) <= temp_mult_18(153);
partial_product_0(154) <= temp_mult_18(154);
partial_product_0(155) <= temp_mult_18(155);
partial_product_0(156) <= temp_mult_18(156);
partial_product_0(157) <= temp_mult_18(157);
partial_product_0(158) <= temp_mult_18(158);
partial_product_0(159) <= temp_mult_18(159);
partial_product_0(160) <= temp_mult_18(160);
partial_product_0(161) <= temp_mult_18(161);
partial_product_0(162) <= temp_mult_18(162);
partial_product_0(163) <= temp_mult_18(163);
partial_product_0(164) <= temp_mult_24(164);
partial_product_0(165) <= temp_mult_24(165);
partial_product_0(166) <= temp_mult_24(166);
partial_product_0(167) <= temp_mult_24(167);
partial_product_0(168) <= temp_mult_24(168);
partial_product_0(169) <= temp_mult_24(169);
partial_product_0(170) <= temp_mult_24(170);
partial_product_0(171) <= temp_mult_24(171);
partial_product_0(172) <= temp_mult_24(172);
partial_product_0(173) <= temp_mult_24(173);
partial_product_0(174) <= temp_mult_24(174);
partial_product_0(175) <= temp_mult_24(175);
partial_product_0(176) <= temp_mult_24(176);
partial_product_0(177) <= temp_mult_24(177);
partial_product_0(178) <= temp_mult_24(178);
partial_product_0(179) <= temp_mult_24(179);
partial_product_0(180) <= temp_mult_24(180);
partial_product_0(181) <= temp_mult_24(181);
partial_product_0(182) <= temp_mult_24(182);
partial_product_0(183) <= temp_mult_24(183);
partial_product_0(184) <= temp_mult_24(184);
partial_product_0(185) <= temp_mult_24(185);
partial_product_0(186) <= temp_mult_24(186);
partial_product_0(187) <= temp_mult_24(187);
partial_product_0(188) <= temp_mult_24(188);
partial_product_0(189) <= temp_mult_24(189);
partial_product_0(190) <= temp_mult_24(190);
partial_product_0(191) <= temp_mult_24(191);
partial_product_0(192) <= temp_mult_24(192);
partial_product_0(193) <= temp_mult_24(193);
partial_product_0(194) <= temp_mult_24(194);
partial_product_0(195) <= temp_mult_24(195);
partial_product_0(196) <= temp_mult_24(196);
partial_product_0(197) <= temp_mult_24(197);
partial_product_0(198) <= temp_mult_24(198);
partial_product_0(199) <= temp_mult_24(199);
partial_product_0(200) <= temp_mult_24(200);
partial_product_0(201) <= temp_mult_24(201);
partial_product_0(202) <= temp_mult_24(202);
partial_product_0(203) <= temp_mult_24(203);
partial_product_0(204) <= temp_mult_24(204);
partial_product_0(205) <= temp_mult_45(205);
partial_product_0(206) <= temp_mult_45(206);
partial_product_0(207) <= temp_mult_45(207);
partial_product_0(208) <= temp_mult_45(208);
partial_product_0(209) <= temp_mult_45(209);
partial_product_0(210) <= temp_mult_45(210);
partial_product_0(211) <= temp_mult_45(211);
partial_product_0(212) <= temp_mult_45(212);
partial_product_0(213) <= temp_mult_45(213);
partial_product_0(214) <= temp_mult_45(214);
partial_product_0(215) <= temp_mult_45(215);
partial_product_0(216) <= temp_mult_45(216);
partial_product_0(217) <= temp_mult_45(217);
partial_product_0(218) <= temp_mult_45(218);
partial_product_0(219) <= temp_mult_45(219);
partial_product_0(220) <= temp_mult_45(220);
partial_product_0(221) <= temp_mult_45(221);
partial_product_0(222) <= temp_mult_45(222);
partial_product_0(223) <= temp_mult_45(223);
partial_product_0(224) <= temp_mult_45(224);
partial_product_0(225) <= temp_mult_45(225);
partial_product_0(226) <= temp_mult_45(226);
partial_product_0(227) <= temp_mult_45(227);
partial_product_0(228) <= temp_mult_45(228);
partial_product_0(229) <= temp_mult_45(229);
partial_product_0(230) <= temp_mult_45(230);
partial_product_0(231) <= temp_mult_45(231);
partial_product_0(232) <= temp_mult_45(232);
partial_product_0(233) <= temp_mult_45(233);
partial_product_0(234) <= temp_mult_45(234);
partial_product_0(235) <= temp_mult_45(235);
partial_product_0(236) <= temp_mult_45(236);
partial_product_0(237) <= temp_mult_45(237);
partial_product_0(238) <= temp_mult_45(238);
partial_product_0(239) <= temp_mult_45(239);
partial_product_0(240) <= temp_mult_45(240);
partial_product_0(241) <= temp_mult_45(241);
partial_product_0(242) <= temp_mult_45(242);
partial_product_0(243) <= temp_mult_45(243);
partial_product_0(244) <= temp_mult_45(244);
partial_product_0(245) <= temp_mult_45(245);
partial_product_0(246) <= temp_mult_54(246);
partial_product_0(247) <= temp_mult_54(247);
partial_product_0(248) <= temp_mult_54(248);
partial_product_0(249) <= temp_mult_54(249);
partial_product_0(250) <= temp_mult_54(250);
partial_product_0(251) <= temp_mult_54(251);
partial_product_0(252) <= temp_mult_54(252);
partial_product_0(253) <= temp_mult_54(253);
partial_product_0(254) <= temp_mult_54(254);
partial_product_0(255) <= temp_mult_54(255);
partial_product_0(256) <= temp_mult_54(256);
partial_product_0(257) <= temp_mult_54(257);
partial_product_0(258) <= temp_mult_54(258);
partial_product_0(259) <= temp_mult_54(259);
partial_product_0(260) <= temp_mult_54(260);
partial_product_0(261) <= temp_mult_54(261);
partial_product_0(262) <= temp_mult_54(262);
partial_product_0(263) <= temp_mult_54(263);
partial_product_0(264) <= temp_mult_54(264);
partial_product_0(265) <= temp_mult_54(265);
partial_product_0(266) <= temp_mult_54(266);
partial_product_0(267) <= temp_mult_54(267);
partial_product_0(268) <= temp_mult_54(268);
partial_product_0(269) <= temp_mult_54(269);
partial_product_0(270) <= temp_mult_54(270);
partial_product_0(271) <= temp_mult_54(271);
partial_product_0(272) <= temp_mult_54(272);
partial_product_0(273) <= temp_mult_54(273);
partial_product_0(274) <= temp_mult_54(274);
partial_product_0(275) <= temp_mult_54(275);
partial_product_0(276) <= temp_mult_54(276);
partial_product_0(277) <= temp_mult_54(277);
partial_product_0(278) <= temp_mult_54(278);
partial_product_0(279) <= temp_mult_54(279);
partial_product_0(280) <= temp_mult_54(280);
partial_product_0(281) <= temp_mult_54(281);
partial_product_0(282) <= temp_mult_54(282);
partial_product_0(283) <= temp_mult_54(283);
partial_product_0(284) <= temp_mult_54(284);
partial_product_0(285) <= temp_mult_54(285);
partial_product_0(286) <= temp_mult_54(286);
partial_product_0(287) <= temp_mult_63(287);
partial_product_0(288) <= temp_mult_63(288);
partial_product_0(289) <= temp_mult_63(289);
partial_product_0(290) <= temp_mult_63(290);
partial_product_0(291) <= temp_mult_63(291);
partial_product_0(292) <= temp_mult_63(292);
partial_product_0(293) <= temp_mult_63(293);
partial_product_0(294) <= temp_mult_63(294);
partial_product_0(295) <= temp_mult_63(295);
partial_product_0(296) <= temp_mult_63(296);
partial_product_0(297) <= temp_mult_63(297);
partial_product_0(298) <= temp_mult_63(298);
partial_product_0(299) <= temp_mult_63(299);
partial_product_0(300) <= temp_mult_63(300);
partial_product_0(301) <= temp_mult_63(301);
partial_product_0(302) <= temp_mult_63(302);
partial_product_0(303) <= temp_mult_63(303);
partial_product_0(304) <= temp_mult_63(304);
partial_product_0(305) <= temp_mult_63(305);
partial_product_0(306) <= temp_mult_63(306);
partial_product_0(307) <= temp_mult_63(307);
partial_product_0(308) <= temp_mult_63(308);
partial_product_0(309) <= temp_mult_63(309);
partial_product_0(310) <= temp_mult_63(310);
partial_product_0(311) <= temp_mult_63(311);
partial_product_0(312) <= temp_mult_63(312);
partial_product_0(313) <= temp_mult_63(313);
partial_product_0(314) <= temp_mult_63(314);
partial_product_0(315) <= temp_mult_63(315);
partial_product_0(316) <= temp_mult_63(316);
partial_product_0(317) <= temp_mult_63(317);
partial_product_0(318) <= temp_mult_63(318);
partial_product_0(319) <= temp_mult_63(319);
partial_product_0(320) <= temp_mult_63(320);
partial_product_0(321) <= temp_mult_63(321);
partial_product_0(322) <= temp_mult_63(322);
partial_product_0(323) <= temp_mult_63(323);
partial_product_0(324) <= temp_mult_63(324);
partial_product_0(325) <= temp_mult_63(325);
partial_product_0(326) <= temp_mult_63(326);
partial_product_0(327) <= temp_mult_63(327);
partial_product_0(328) <= temp_mult_123(328);
partial_product_0(329) <= temp_mult_123(329);
partial_product_0(330) <= temp_mult_123(330);
partial_product_0(331) <= temp_mult_123(331);
partial_product_0(332) <= temp_mult_123(332);
partial_product_0(333) <= temp_mult_123(333);
partial_product_0(334) <= temp_mult_123(334);
partial_product_0(335) <= temp_mult_123(335);
partial_product_0(336) <= temp_mult_123(336);
partial_product_0(337) <= temp_mult_123(337);
partial_product_0(338) <= temp_mult_123(338);
partial_product_0(339) <= temp_mult_123(339);
partial_product_0(340) <= temp_mult_123(340);
partial_product_0(341) <= temp_mult_123(341);
partial_product_0(342) <= temp_mult_123(342);
partial_product_0(343) <= temp_mult_123(343);
partial_product_0(344) <= temp_mult_123(344);
partial_product_0(345) <= temp_mult_123(345);
partial_product_0(346) <= temp_mult_123(346);
partial_product_0(347) <= temp_mult_123(347);
partial_product_0(348) <= temp_mult_123(348);
partial_product_0(349) <= temp_mult_123(349);
partial_product_0(350) <= temp_mult_123(350);
partial_product_0(351) <= temp_mult_123(351);
partial_product_0(352) <= temp_mult_123(352);
partial_product_0(353) <= temp_mult_123(353);
partial_product_0(354) <= temp_mult_123(354);
partial_product_0(355) <= temp_mult_123(355);
partial_product_0(356) <= temp_mult_123(356);
partial_product_0(357) <= temp_mult_123(357);
partial_product_0(358) <= temp_mult_123(358);
partial_product_0(359) <= temp_mult_123(359);
partial_product_0(360) <= temp_mult_123(360);
partial_product_0(361) <= temp_mult_123(361);
partial_product_0(362) <= temp_mult_123(362);
partial_product_0(363) <= temp_mult_123(363);
partial_product_0(364) <= temp_mult_123(364);
partial_product_0(365) <= temp_mult_123(365);
partial_product_0(366) <= temp_mult_123(366);
partial_product_0(367) <= temp_mult_123(367);
partial_product_0(368) <= temp_mult_123(368);
partial_product_0(369) <= temp_mult_129(369);
partial_product_0(370) <= temp_mult_129(370);
partial_product_0(371) <= temp_mult_129(371);
partial_product_0(372) <= temp_mult_129(372);
partial_product_0(373) <= temp_mult_129(373);
partial_product_0(374) <= temp_mult_129(374);
partial_product_0(375) <= temp_mult_129(375);
partial_product_0(376) <= temp_mult_129(376);
partial_product_0(377) <= temp_mult_129(377);
partial_product_0(378) <= temp_mult_129(378);
partial_product_0(379) <= temp_mult_129(379);
partial_product_0(380) <= temp_mult_129(380);
partial_product_0(381) <= temp_mult_129(381);
partial_product_0(382) <= temp_mult_129(382);
partial_product_0(383) <= temp_mult_129(383);
partial_product_0(384) <= temp_mult_129(384);
partial_product_0(385) <= temp_mult_129(385);
partial_product_0(386) <= temp_mult_129(386);
partial_product_0(387) <= temp_mult_129(387);
partial_product_0(388) <= temp_mult_129(388);
partial_product_0(389) <= temp_mult_129(389);
partial_product_0(390) <= temp_mult_129(390);
partial_product_0(391) <= temp_mult_129(391);
partial_product_0(392) <= temp_mult_129(392);
partial_product_0(393) <= temp_mult_129(393);
partial_product_0(394) <= temp_mult_129(394);
partial_product_0(395) <= temp_mult_129(395);
partial_product_0(396) <= temp_mult_129(396);
partial_product_0(397) <= temp_mult_129(397);
partial_product_0(398) <= temp_mult_129(398);
partial_product_0(399) <= temp_mult_129(399);
partial_product_0(400) <= temp_mult_129(400);
partial_product_0(401) <= temp_mult_129(401);
partial_product_0(402) <= temp_mult_129(402);
partial_product_0(403) <= temp_mult_129(403);
partial_product_0(404) <= temp_mult_129(404);
partial_product_0(405) <= temp_mult_129(405);
partial_product_0(406) <= temp_mult_129(406);
partial_product_0(407) <= temp_mult_129(407);
partial_product_0(408) <= temp_mult_129(408);
partial_product_0(409) <= temp_mult_129(409);
partial_product_0(410) <= '0';
partial_product_0(411) <= '0';
partial_product_0(412) <= '0';
partial_product_0(413) <= temp_mult_148(413);
partial_product_0(414) <= temp_mult_148(414);
partial_product_0(415) <= temp_mult_148(415);
partial_product_0(416) <= temp_mult_148(416);
partial_product_0(417) <= temp_mult_148(417);
partial_product_0(418) <= temp_mult_148(418);
partial_product_0(419) <= temp_mult_148(419);
partial_product_0(420) <= temp_mult_148(420);
partial_product_0(421) <= temp_mult_148(421);
partial_product_0(422) <= temp_mult_148(422);
partial_product_0(423) <= temp_mult_148(423);
partial_product_0(424) <= temp_mult_148(424);
partial_product_0(425) <= temp_mult_148(425);
partial_product_0(426) <= temp_mult_148(426);
partial_product_0(427) <= temp_mult_148(427);
partial_product_0(428) <= temp_mult_148(428);
partial_product_0(429) <= temp_mult_148(429);
partial_product_0(430) <= temp_mult_148(430);
partial_product_0(431) <= temp_mult_148(431);
partial_product_0(432) <= temp_mult_148(432);
partial_product_0(433) <= temp_mult_148(433);
partial_product_0(434) <= temp_mult_148(434);
partial_product_0(435) <= temp_mult_148(435);
partial_product_0(436) <= temp_mult_148(436);
partial_product_0(437) <= temp_mult_148(437);
partial_product_0(438) <= temp_mult_148(438);
partial_product_0(439) <= temp_mult_148(439);
partial_product_0(440) <= temp_mult_148(440);
partial_product_0(441) <= temp_mult_148(441);
partial_product_0(442) <= temp_mult_148(442);
partial_product_0(443) <= temp_mult_148(443);
partial_product_0(444) <= temp_mult_148(444);
partial_product_0(445) <= temp_mult_148(445);
partial_product_0(446) <= temp_mult_148(446);
partial_product_0(447) <= temp_mult_148(447);
partial_product_0(448) <= temp_mult_148(448);
partial_product_0(449) <= temp_mult_148(449);
partial_product_0(450) <= temp_mult_148(450);
partial_product_0(451) <= temp_mult_148(451);
partial_product_0(452) <= temp_mult_148(452);
partial_product_0(453) <= temp_mult_148(453);
partial_product_0(454) <= temp_mult_154(454);
partial_product_0(455) <= temp_mult_154(455);
partial_product_0(456) <= temp_mult_154(456);
partial_product_0(457) <= temp_mult_154(457);
partial_product_0(458) <= temp_mult_154(458);
partial_product_0(459) <= temp_mult_154(459);
partial_product_0(460) <= temp_mult_154(460);
partial_product_0(461) <= temp_mult_154(461);
partial_product_0(462) <= temp_mult_154(462);
partial_product_0(463) <= temp_mult_154(463);
partial_product_0(464) <= temp_mult_154(464);
partial_product_0(465) <= temp_mult_154(465);
partial_product_0(466) <= temp_mult_154(466);
partial_product_0(467) <= temp_mult_154(467);
partial_product_0(468) <= temp_mult_154(468);
partial_product_0(469) <= temp_mult_154(469);
partial_product_0(470) <= temp_mult_154(470);
partial_product_0(471) <= temp_mult_154(471);
partial_product_0(472) <= temp_mult_154(472);
partial_product_0(473) <= temp_mult_154(473);
partial_product_0(474) <= temp_mult_154(474);
partial_product_0(475) <= temp_mult_154(475);
partial_product_0(476) <= temp_mult_154(476);
partial_product_0(477) <= temp_mult_154(477);
partial_product_0(478) <= temp_mult_154(478);
partial_product_0(479) <= temp_mult_154(479);
partial_product_0(480) <= temp_mult_154(480);
partial_product_0(481) <= temp_mult_154(481);
partial_product_0(482) <= temp_mult_154(482);
partial_product_0(483) <= temp_mult_154(483);
partial_product_0(484) <= temp_mult_154(484);
partial_product_0(485) <= temp_mult_154(485);
partial_product_0(486) <= temp_mult_154(486);
partial_product_0(487) <= temp_mult_154(487);
partial_product_0(488) <= temp_mult_154(488);
partial_product_0(489) <= temp_mult_154(489);
partial_product_0(490) <= temp_mult_154(490);
partial_product_0(491) <= temp_mult_154(491);
partial_product_0(492) <= temp_mult_154(492);
partial_product_0(493) <= temp_mult_154(493);
partial_product_0(494) <= temp_mult_154(494);
partial_product_0(495) <= '0';
partial_product_0(496) <= '0';
partial_product_0(497) <= '0';
partial_product_0(498) <= '0';
partial_product_0(499) <= '0';
partial_product_0(500) <= '0';
partial_product_0(501) <= '0';
partial_product_0(502) <= '0';
partial_product_0(503) <= '0';
partial_product_0(504) <= '0';
partial_product_0(505) <= '0';
partial_product_0(506) <= '0';
partial_product_0(507) <= '0';
partial_product_0(508) <= '0';
partial_product_0(509) <= '0';
partial_product_0(510) <= '0';
partial_product_0(511) <= '0';
partial_product_0(512) <= '0';
partial_product_1(0) <= '0';
partial_product_1(1) <= '0';
partial_product_1(2) <= '0';
partial_product_1(3) <= '0';
partial_product_1(4) <= '0';
partial_product_1(5) <= '0';
partial_product_1(6) <= '0';
partial_product_1(7) <= '0';
partial_product_1(8) <= '0';
partial_product_1(9) <= '0';
partial_product_1(10) <= '0';
partial_product_1(11) <= '0';
partial_product_1(12) <= '0';
partial_product_1(13) <= '0';
partial_product_1(14) <= '0';
partial_product_1(15) <= '0';
partial_product_1(16) <= '0';
partial_product_1(17) <= temp_mult_5(17);
partial_product_1(18) <= temp_mult_5(18);
partial_product_1(19) <= temp_mult_5(19);
partial_product_1(20) <= temp_mult_5(20);
partial_product_1(21) <= temp_mult_5(21);
partial_product_1(22) <= temp_mult_5(22);
partial_product_1(23) <= temp_mult_5(23);
partial_product_1(24) <= temp_mult_5(24);
partial_product_1(25) <= temp_mult_5(25);
partial_product_1(26) <= temp_mult_5(26);
partial_product_1(27) <= temp_mult_5(27);
partial_product_1(28) <= temp_mult_5(28);
partial_product_1(29) <= temp_mult_5(29);
partial_product_1(30) <= temp_mult_5(30);
partial_product_1(31) <= temp_mult_5(31);
partial_product_1(32) <= temp_mult_5(32);
partial_product_1(33) <= temp_mult_5(33);
partial_product_1(34) <= temp_mult_5(34);
partial_product_1(35) <= temp_mult_5(35);
partial_product_1(36) <= temp_mult_5(36);
partial_product_1(37) <= temp_mult_5(37);
partial_product_1(38) <= temp_mult_5(38);
partial_product_1(39) <= temp_mult_5(39);
partial_product_1(40) <= temp_mult_5(40);
partial_product_1(41) <= temp_mult_5(41);
partial_product_1(42) <= temp_mult_5(42);
partial_product_1(43) <= temp_mult_5(43);
partial_product_1(44) <= temp_mult_5(44);
partial_product_1(45) <= temp_mult_5(45);
partial_product_1(46) <= temp_mult_5(46);
partial_product_1(47) <= temp_mult_5(47);
partial_product_1(48) <= temp_mult_5(48);
partial_product_1(49) <= temp_mult_5(49);
partial_product_1(50) <= temp_mult_5(50);
partial_product_1(51) <= temp_mult_5(51);
partial_product_1(52) <= temp_mult_5(52);
partial_product_1(53) <= temp_mult_5(53);
partial_product_1(54) <= temp_mult_5(54);
partial_product_1(55) <= temp_mult_5(55);
partial_product_1(56) <= temp_mult_5(56);
partial_product_1(57) <= temp_mult_5(57);
partial_product_1(58) <= temp_mult_11(58);
partial_product_1(59) <= temp_mult_11(59);
partial_product_1(60) <= temp_mult_11(60);
partial_product_1(61) <= temp_mult_11(61);
partial_product_1(62) <= temp_mult_11(62);
partial_product_1(63) <= temp_mult_11(63);
partial_product_1(64) <= temp_mult_11(64);
partial_product_1(65) <= temp_mult_11(65);
partial_product_1(66) <= temp_mult_11(66);
partial_product_1(67) <= temp_mult_11(67);
partial_product_1(68) <= temp_mult_11(68);
partial_product_1(69) <= temp_mult_11(69);
partial_product_1(70) <= temp_mult_11(70);
partial_product_1(71) <= temp_mult_11(71);
partial_product_1(72) <= temp_mult_11(72);
partial_product_1(73) <= temp_mult_11(73);
partial_product_1(74) <= temp_mult_11(74);
partial_product_1(75) <= temp_mult_11(75);
partial_product_1(76) <= temp_mult_11(76);
partial_product_1(77) <= temp_mult_11(77);
partial_product_1(78) <= temp_mult_11(78);
partial_product_1(79) <= temp_mult_11(79);
partial_product_1(80) <= temp_mult_11(80);
partial_product_1(81) <= temp_mult_11(81);
partial_product_1(82) <= temp_mult_11(82);
partial_product_1(83) <= temp_mult_11(83);
partial_product_1(84) <= temp_mult_11(84);
partial_product_1(85) <= temp_mult_11(85);
partial_product_1(86) <= temp_mult_11(86);
partial_product_1(87) <= temp_mult_11(87);
partial_product_1(88) <= temp_mult_11(88);
partial_product_1(89) <= temp_mult_11(89);
partial_product_1(90) <= temp_mult_11(90);
partial_product_1(91) <= temp_mult_11(91);
partial_product_1(92) <= temp_mult_11(92);
partial_product_1(93) <= temp_mult_11(93);
partial_product_1(94) <= temp_mult_11(94);
partial_product_1(95) <= temp_mult_11(95);
partial_product_1(96) <= temp_mult_11(96);
partial_product_1(97) <= temp_mult_11(97);
partial_product_1(98) <= temp_mult_11(98);
partial_product_1(99) <= temp_mult_17(99);
partial_product_1(100) <= temp_mult_17(100);
partial_product_1(101) <= temp_mult_17(101);
partial_product_1(102) <= temp_mult_17(102);
partial_product_1(103) <= temp_mult_17(103);
partial_product_1(104) <= temp_mult_17(104);
partial_product_1(105) <= temp_mult_17(105);
partial_product_1(106) <= temp_mult_17(106);
partial_product_1(107) <= temp_mult_17(107);
partial_product_1(108) <= temp_mult_17(108);
partial_product_1(109) <= temp_mult_17(109);
partial_product_1(110) <= temp_mult_17(110);
partial_product_1(111) <= temp_mult_17(111);
partial_product_1(112) <= temp_mult_17(112);
partial_product_1(113) <= temp_mult_17(113);
partial_product_1(114) <= temp_mult_17(114);
partial_product_1(115) <= temp_mult_17(115);
partial_product_1(116) <= temp_mult_17(116);
partial_product_1(117) <= temp_mult_17(117);
partial_product_1(118) <= temp_mult_17(118);
partial_product_1(119) <= temp_mult_17(119);
partial_product_1(120) <= temp_mult_17(120);
partial_product_1(121) <= temp_mult_17(121);
partial_product_1(122) <= temp_mult_17(122);
partial_product_1(123) <= temp_mult_17(123);
partial_product_1(124) <= temp_mult_17(124);
partial_product_1(125) <= temp_mult_17(125);
partial_product_1(126) <= temp_mult_17(126);
partial_product_1(127) <= temp_mult_17(127);
partial_product_1(128) <= temp_mult_17(128);
partial_product_1(129) <= temp_mult_17(129);
partial_product_1(130) <= temp_mult_17(130);
partial_product_1(131) <= temp_mult_17(131);
partial_product_1(132) <= temp_mult_17(132);
partial_product_1(133) <= temp_mult_17(133);
partial_product_1(134) <= temp_mult_17(134);
partial_product_1(135) <= temp_mult_17(135);
partial_product_1(136) <= temp_mult_17(136);
partial_product_1(137) <= temp_mult_17(137);
partial_product_1(138) <= temp_mult_17(138);
partial_product_1(139) <= temp_mult_17(139);
partial_product_1(140) <= temp_mult_23(140);
partial_product_1(141) <= temp_mult_23(141);
partial_product_1(142) <= temp_mult_23(142);
partial_product_1(143) <= temp_mult_23(143);
partial_product_1(144) <= temp_mult_23(144);
partial_product_1(145) <= temp_mult_23(145);
partial_product_1(146) <= temp_mult_23(146);
partial_product_1(147) <= temp_mult_23(147);
partial_product_1(148) <= temp_mult_23(148);
partial_product_1(149) <= temp_mult_23(149);
partial_product_1(150) <= temp_mult_23(150);
partial_product_1(151) <= temp_mult_23(151);
partial_product_1(152) <= temp_mult_23(152);
partial_product_1(153) <= temp_mult_23(153);
partial_product_1(154) <= temp_mult_23(154);
partial_product_1(155) <= temp_mult_23(155);
partial_product_1(156) <= temp_mult_23(156);
partial_product_1(157) <= temp_mult_23(157);
partial_product_1(158) <= temp_mult_23(158);
partial_product_1(159) <= temp_mult_23(159);
partial_product_1(160) <= temp_mult_23(160);
partial_product_1(161) <= temp_mult_23(161);
partial_product_1(162) <= temp_mult_23(162);
partial_product_1(163) <= temp_mult_23(163);
partial_product_1(164) <= temp_mult_23(164);
partial_product_1(165) <= temp_mult_23(165);
partial_product_1(166) <= temp_mult_23(166);
partial_product_1(167) <= temp_mult_23(167);
partial_product_1(168) <= temp_mult_23(168);
partial_product_1(169) <= temp_mult_23(169);
partial_product_1(170) <= temp_mult_23(170);
partial_product_1(171) <= temp_mult_23(171);
partial_product_1(172) <= temp_mult_23(172);
partial_product_1(173) <= temp_mult_23(173);
partial_product_1(174) <= temp_mult_23(174);
partial_product_1(175) <= temp_mult_23(175);
partial_product_1(176) <= temp_mult_23(176);
partial_product_1(177) <= temp_mult_23(177);
partial_product_1(178) <= temp_mult_23(178);
partial_product_1(179) <= temp_mult_23(179);
partial_product_1(180) <= temp_mult_23(180);
partial_product_1(181) <= temp_mult_29(181);
partial_product_1(182) <= temp_mult_29(182);
partial_product_1(183) <= temp_mult_29(183);
partial_product_1(184) <= temp_mult_29(184);
partial_product_1(185) <= temp_mult_29(185);
partial_product_1(186) <= temp_mult_29(186);
partial_product_1(187) <= temp_mult_29(187);
partial_product_1(188) <= temp_mult_29(188);
partial_product_1(189) <= temp_mult_29(189);
partial_product_1(190) <= temp_mult_29(190);
partial_product_1(191) <= temp_mult_29(191);
partial_product_1(192) <= temp_mult_29(192);
partial_product_1(193) <= temp_mult_29(193);
partial_product_1(194) <= temp_mult_29(194);
partial_product_1(195) <= temp_mult_29(195);
partial_product_1(196) <= temp_mult_29(196);
partial_product_1(197) <= temp_mult_29(197);
partial_product_1(198) <= temp_mult_29(198);
partial_product_1(199) <= temp_mult_29(199);
partial_product_1(200) <= temp_mult_29(200);
partial_product_1(201) <= temp_mult_29(201);
partial_product_1(202) <= temp_mult_29(202);
partial_product_1(203) <= temp_mult_29(203);
partial_product_1(204) <= temp_mult_29(204);
partial_product_1(205) <= temp_mult_29(205);
partial_product_1(206) <= temp_mult_29(206);
partial_product_1(207) <= temp_mult_29(207);
partial_product_1(208) <= temp_mult_29(208);
partial_product_1(209) <= temp_mult_29(209);
partial_product_1(210) <= temp_mult_29(210);
partial_product_1(211) <= temp_mult_29(211);
partial_product_1(212) <= temp_mult_29(212);
partial_product_1(213) <= temp_mult_29(213);
partial_product_1(214) <= temp_mult_29(214);
partial_product_1(215) <= temp_mult_29(215);
partial_product_1(216) <= temp_mult_29(216);
partial_product_1(217) <= temp_mult_29(217);
partial_product_1(218) <= temp_mult_29(218);
partial_product_1(219) <= temp_mult_29(219);
partial_product_1(220) <= temp_mult_29(220);
partial_product_1(221) <= temp_mult_29(221);
partial_product_1(222) <= temp_mult_46(222);
partial_product_1(223) <= temp_mult_46(223);
partial_product_1(224) <= temp_mult_46(224);
partial_product_1(225) <= temp_mult_46(225);
partial_product_1(226) <= temp_mult_46(226);
partial_product_1(227) <= temp_mult_46(227);
partial_product_1(228) <= temp_mult_46(228);
partial_product_1(229) <= temp_mult_46(229);
partial_product_1(230) <= temp_mult_46(230);
partial_product_1(231) <= temp_mult_46(231);
partial_product_1(232) <= temp_mult_46(232);
partial_product_1(233) <= temp_mult_46(233);
partial_product_1(234) <= temp_mult_46(234);
partial_product_1(235) <= temp_mult_46(235);
partial_product_1(236) <= temp_mult_46(236);
partial_product_1(237) <= temp_mult_46(237);
partial_product_1(238) <= temp_mult_46(238);
partial_product_1(239) <= temp_mult_46(239);
partial_product_1(240) <= temp_mult_46(240);
partial_product_1(241) <= temp_mult_46(241);
partial_product_1(242) <= temp_mult_46(242);
partial_product_1(243) <= temp_mult_46(243);
partial_product_1(244) <= temp_mult_46(244);
partial_product_1(245) <= temp_mult_46(245);
partial_product_1(246) <= temp_mult_46(246);
partial_product_1(247) <= temp_mult_46(247);
partial_product_1(248) <= temp_mult_46(248);
partial_product_1(249) <= temp_mult_46(249);
partial_product_1(250) <= temp_mult_46(250);
partial_product_1(251) <= temp_mult_46(251);
partial_product_1(252) <= temp_mult_46(252);
partial_product_1(253) <= temp_mult_46(253);
partial_product_1(254) <= temp_mult_46(254);
partial_product_1(255) <= temp_mult_46(255);
partial_product_1(256) <= temp_mult_46(256);
partial_product_1(257) <= temp_mult_46(257);
partial_product_1(258) <= temp_mult_46(258);
partial_product_1(259) <= temp_mult_46(259);
partial_product_1(260) <= temp_mult_46(260);
partial_product_1(261) <= temp_mult_46(261);
partial_product_1(262) <= temp_mult_46(262);
partial_product_1(263) <= temp_mult_55(263);
partial_product_1(264) <= temp_mult_55(264);
partial_product_1(265) <= temp_mult_55(265);
partial_product_1(266) <= temp_mult_55(266);
partial_product_1(267) <= temp_mult_55(267);
partial_product_1(268) <= temp_mult_55(268);
partial_product_1(269) <= temp_mult_55(269);
partial_product_1(270) <= temp_mult_55(270);
partial_product_1(271) <= temp_mult_55(271);
partial_product_1(272) <= temp_mult_55(272);
partial_product_1(273) <= temp_mult_55(273);
partial_product_1(274) <= temp_mult_55(274);
partial_product_1(275) <= temp_mult_55(275);
partial_product_1(276) <= temp_mult_55(276);
partial_product_1(277) <= temp_mult_55(277);
partial_product_1(278) <= temp_mult_55(278);
partial_product_1(279) <= temp_mult_55(279);
partial_product_1(280) <= temp_mult_55(280);
partial_product_1(281) <= temp_mult_55(281);
partial_product_1(282) <= temp_mult_55(282);
partial_product_1(283) <= temp_mult_55(283);
partial_product_1(284) <= temp_mult_55(284);
partial_product_1(285) <= temp_mult_55(285);
partial_product_1(286) <= temp_mult_55(286);
partial_product_1(287) <= temp_mult_55(287);
partial_product_1(288) <= temp_mult_55(288);
partial_product_1(289) <= temp_mult_55(289);
partial_product_1(290) <= temp_mult_55(290);
partial_product_1(291) <= temp_mult_55(291);
partial_product_1(292) <= temp_mult_55(292);
partial_product_1(293) <= temp_mult_55(293);
partial_product_1(294) <= temp_mult_55(294);
partial_product_1(295) <= temp_mult_55(295);
partial_product_1(296) <= temp_mult_55(296);
partial_product_1(297) <= temp_mult_55(297);
partial_product_1(298) <= temp_mult_55(298);
partial_product_1(299) <= temp_mult_55(299);
partial_product_1(300) <= temp_mult_55(300);
partial_product_1(301) <= temp_mult_55(301);
partial_product_1(302) <= temp_mult_55(302);
partial_product_1(303) <= temp_mult_55(303);
partial_product_1(304) <= temp_mult_122(304);
partial_product_1(305) <= temp_mult_122(305);
partial_product_1(306) <= temp_mult_122(306);
partial_product_1(307) <= temp_mult_122(307);
partial_product_1(308) <= temp_mult_122(308);
partial_product_1(309) <= temp_mult_122(309);
partial_product_1(310) <= temp_mult_122(310);
partial_product_1(311) <= temp_mult_122(311);
partial_product_1(312) <= temp_mult_122(312);
partial_product_1(313) <= temp_mult_122(313);
partial_product_1(314) <= temp_mult_122(314);
partial_product_1(315) <= temp_mult_122(315);
partial_product_1(316) <= temp_mult_122(316);
partial_product_1(317) <= temp_mult_122(317);
partial_product_1(318) <= temp_mult_122(318);
partial_product_1(319) <= temp_mult_122(319);
partial_product_1(320) <= temp_mult_122(320);
partial_product_1(321) <= temp_mult_122(321);
partial_product_1(322) <= temp_mult_122(322);
partial_product_1(323) <= temp_mult_122(323);
partial_product_1(324) <= temp_mult_122(324);
partial_product_1(325) <= temp_mult_122(325);
partial_product_1(326) <= temp_mult_122(326);
partial_product_1(327) <= temp_mult_122(327);
partial_product_1(328) <= temp_mult_122(328);
partial_product_1(329) <= temp_mult_122(329);
partial_product_1(330) <= temp_mult_122(330);
partial_product_1(331) <= temp_mult_122(331);
partial_product_1(332) <= temp_mult_122(332);
partial_product_1(333) <= temp_mult_122(333);
partial_product_1(334) <= temp_mult_122(334);
partial_product_1(335) <= temp_mult_122(335);
partial_product_1(336) <= temp_mult_122(336);
partial_product_1(337) <= temp_mult_122(337);
partial_product_1(338) <= temp_mult_122(338);
partial_product_1(339) <= temp_mult_122(339);
partial_product_1(340) <= temp_mult_122(340);
partial_product_1(341) <= temp_mult_122(341);
partial_product_1(342) <= temp_mult_122(342);
partial_product_1(343) <= temp_mult_122(343);
partial_product_1(344) <= temp_mult_122(344);
partial_product_1(345) <= temp_mult_128(345);
partial_product_1(346) <= temp_mult_128(346);
partial_product_1(347) <= temp_mult_128(347);
partial_product_1(348) <= temp_mult_128(348);
partial_product_1(349) <= temp_mult_128(349);
partial_product_1(350) <= temp_mult_128(350);
partial_product_1(351) <= temp_mult_128(351);
partial_product_1(352) <= temp_mult_128(352);
partial_product_1(353) <= temp_mult_128(353);
partial_product_1(354) <= temp_mult_128(354);
partial_product_1(355) <= temp_mult_128(355);
partial_product_1(356) <= temp_mult_128(356);
partial_product_1(357) <= temp_mult_128(357);
partial_product_1(358) <= temp_mult_128(358);
partial_product_1(359) <= temp_mult_128(359);
partial_product_1(360) <= temp_mult_128(360);
partial_product_1(361) <= temp_mult_128(361);
partial_product_1(362) <= temp_mult_128(362);
partial_product_1(363) <= temp_mult_128(363);
partial_product_1(364) <= temp_mult_128(364);
partial_product_1(365) <= temp_mult_128(365);
partial_product_1(366) <= temp_mult_128(366);
partial_product_1(367) <= temp_mult_128(367);
partial_product_1(368) <= temp_mult_128(368);
partial_product_1(369) <= temp_mult_128(369);
partial_product_1(370) <= temp_mult_128(370);
partial_product_1(371) <= temp_mult_128(371);
partial_product_1(372) <= temp_mult_128(372);
partial_product_1(373) <= temp_mult_128(373);
partial_product_1(374) <= temp_mult_128(374);
partial_product_1(375) <= temp_mult_128(375);
partial_product_1(376) <= temp_mult_128(376);
partial_product_1(377) <= temp_mult_128(377);
partial_product_1(378) <= temp_mult_128(378);
partial_product_1(379) <= temp_mult_128(379);
partial_product_1(380) <= temp_mult_128(380);
partial_product_1(381) <= temp_mult_128(381);
partial_product_1(382) <= temp_mult_128(382);
partial_product_1(383) <= temp_mult_128(383);
partial_product_1(384) <= temp_mult_128(384);
partial_product_1(385) <= temp_mult_128(385);
partial_product_1(386) <= temp_mult_134(386);
partial_product_1(387) <= temp_mult_134(387);
partial_product_1(388) <= temp_mult_134(388);
partial_product_1(389) <= temp_mult_134(389);
partial_product_1(390) <= temp_mult_134(390);
partial_product_1(391) <= temp_mult_134(391);
partial_product_1(392) <= temp_mult_134(392);
partial_product_1(393) <= temp_mult_134(393);
partial_product_1(394) <= temp_mult_134(394);
partial_product_1(395) <= temp_mult_134(395);
partial_product_1(396) <= temp_mult_134(396);
partial_product_1(397) <= temp_mult_134(397);
partial_product_1(398) <= temp_mult_134(398);
partial_product_1(399) <= temp_mult_134(399);
partial_product_1(400) <= temp_mult_134(400);
partial_product_1(401) <= temp_mult_134(401);
partial_product_1(402) <= temp_mult_134(402);
partial_product_1(403) <= temp_mult_134(403);
partial_product_1(404) <= temp_mult_134(404);
partial_product_1(405) <= temp_mult_134(405);
partial_product_1(406) <= temp_mult_134(406);
partial_product_1(407) <= temp_mult_134(407);
partial_product_1(408) <= temp_mult_134(408);
partial_product_1(409) <= temp_mult_134(409);
partial_product_1(410) <= temp_mult_134(410);
partial_product_1(411) <= temp_mult_134(411);
partial_product_1(412) <= temp_mult_134(412);
partial_product_1(413) <= temp_mult_134(413);
partial_product_1(414) <= temp_mult_134(414);
partial_product_1(415) <= temp_mult_134(415);
partial_product_1(416) <= temp_mult_134(416);
partial_product_1(417) <= temp_mult_134(417);
partial_product_1(418) <= temp_mult_134(418);
partial_product_1(419) <= temp_mult_134(419);
partial_product_1(420) <= temp_mult_134(420);
partial_product_1(421) <= temp_mult_134(421);
partial_product_1(422) <= temp_mult_134(422);
partial_product_1(423) <= temp_mult_134(423);
partial_product_1(424) <= temp_mult_134(424);
partial_product_1(425) <= temp_mult_134(425);
partial_product_1(426) <= temp_mult_134(426);
partial_product_1(427) <= '0';
partial_product_1(428) <= '0';
partial_product_1(429) <= '0';
partial_product_1(430) <= temp_mult_153(430);
partial_product_1(431) <= temp_mult_153(431);
partial_product_1(432) <= temp_mult_153(432);
partial_product_1(433) <= temp_mult_153(433);
partial_product_1(434) <= temp_mult_153(434);
partial_product_1(435) <= temp_mult_153(435);
partial_product_1(436) <= temp_mult_153(436);
partial_product_1(437) <= temp_mult_153(437);
partial_product_1(438) <= temp_mult_153(438);
partial_product_1(439) <= temp_mult_153(439);
partial_product_1(440) <= temp_mult_153(440);
partial_product_1(441) <= temp_mult_153(441);
partial_product_1(442) <= temp_mult_153(442);
partial_product_1(443) <= temp_mult_153(443);
partial_product_1(444) <= temp_mult_153(444);
partial_product_1(445) <= temp_mult_153(445);
partial_product_1(446) <= temp_mult_153(446);
partial_product_1(447) <= temp_mult_153(447);
partial_product_1(448) <= temp_mult_153(448);
partial_product_1(449) <= temp_mult_153(449);
partial_product_1(450) <= temp_mult_153(450);
partial_product_1(451) <= temp_mult_153(451);
partial_product_1(452) <= temp_mult_153(452);
partial_product_1(453) <= temp_mult_153(453);
partial_product_1(454) <= temp_mult_153(454);
partial_product_1(455) <= temp_mult_153(455);
partial_product_1(456) <= temp_mult_153(456);
partial_product_1(457) <= temp_mult_153(457);
partial_product_1(458) <= temp_mult_153(458);
partial_product_1(459) <= temp_mult_153(459);
partial_product_1(460) <= temp_mult_153(460);
partial_product_1(461) <= temp_mult_153(461);
partial_product_1(462) <= temp_mult_153(462);
partial_product_1(463) <= temp_mult_153(463);
partial_product_1(464) <= temp_mult_153(464);
partial_product_1(465) <= temp_mult_153(465);
partial_product_1(466) <= temp_mult_153(466);
partial_product_1(467) <= temp_mult_153(467);
partial_product_1(468) <= temp_mult_153(468);
partial_product_1(469) <= temp_mult_153(469);
partial_product_1(470) <= temp_mult_153(470);
partial_product_1(471) <= temp_mult_159(471);
partial_product_1(472) <= temp_mult_159(472);
partial_product_1(473) <= temp_mult_159(473);
partial_product_1(474) <= temp_mult_159(474);
partial_product_1(475) <= temp_mult_159(475);
partial_product_1(476) <= temp_mult_159(476);
partial_product_1(477) <= temp_mult_159(477);
partial_product_1(478) <= temp_mult_159(478);
partial_product_1(479) <= temp_mult_159(479);
partial_product_1(480) <= temp_mult_159(480);
partial_product_1(481) <= temp_mult_159(481);
partial_product_1(482) <= temp_mult_159(482);
partial_product_1(483) <= temp_mult_159(483);
partial_product_1(484) <= temp_mult_159(484);
partial_product_1(485) <= temp_mult_159(485);
partial_product_1(486) <= temp_mult_159(486);
partial_product_1(487) <= temp_mult_159(487);
partial_product_1(488) <= temp_mult_159(488);
partial_product_1(489) <= temp_mult_159(489);
partial_product_1(490) <= temp_mult_159(490);
partial_product_1(491) <= temp_mult_159(491);
partial_product_1(492) <= temp_mult_159(492);
partial_product_1(493) <= temp_mult_159(493);
partial_product_1(494) <= temp_mult_159(494);
partial_product_1(495) <= temp_mult_159(495);
partial_product_1(496) <= temp_mult_159(496);
partial_product_1(497) <= temp_mult_159(497);
partial_product_1(498) <= temp_mult_159(498);
partial_product_1(499) <= temp_mult_159(499);
partial_product_1(500) <= temp_mult_159(500);
partial_product_1(501) <= temp_mult_159(501);
partial_product_1(502) <= temp_mult_159(502);
partial_product_1(503) <= temp_mult_159(503);
partial_product_1(504) <= temp_mult_159(504);
partial_product_1(505) <= temp_mult_159(505);
partial_product_1(506) <= temp_mult_159(506);
partial_product_1(507) <= temp_mult_159(507);
partial_product_1(508) <= temp_mult_159(508);
partial_product_1(509) <= temp_mult_159(509);
partial_product_1(510) <= temp_mult_159(510);
partial_product_1(511) <= temp_mult_159(511);
partial_product_1(512) <= '0';
partial_product_2(0) <= '0';
partial_product_2(1) <= '0';
partial_product_2(2) <= '0';
partial_product_2(3) <= '0';
partial_product_2(4) <= '0';
partial_product_2(5) <= '0';
partial_product_2(6) <= '0';
partial_product_2(7) <= '0';
partial_product_2(8) <= '0';
partial_product_2(9) <= '0';
partial_product_2(10) <= '0';
partial_product_2(11) <= '0';
partial_product_2(12) <= '0';
partial_product_2(13) <= '0';
partial_product_2(14) <= '0';
partial_product_2(15) <= '0';
partial_product_2(16) <= '0';
partial_product_2(17) <= '0';
partial_product_2(18) <= '0';
partial_product_2(19) <= '0';
partial_product_2(20) <= '0';
partial_product_2(21) <= '0';
partial_product_2(22) <= '0';
partial_product_2(23) <= '0';
partial_product_2(24) <= temp_mult_1(24);
partial_product_2(25) <= temp_mult_1(25);
partial_product_2(26) <= temp_mult_1(26);
partial_product_2(27) <= temp_mult_1(27);
partial_product_2(28) <= temp_mult_1(28);
partial_product_2(29) <= temp_mult_1(29);
partial_product_2(30) <= temp_mult_1(30);
partial_product_2(31) <= temp_mult_1(31);
partial_product_2(32) <= temp_mult_1(32);
partial_product_2(33) <= temp_mult_1(33);
partial_product_2(34) <= temp_mult_1(34);
partial_product_2(35) <= temp_mult_1(35);
partial_product_2(36) <= temp_mult_1(36);
partial_product_2(37) <= temp_mult_1(37);
partial_product_2(38) <= temp_mult_1(38);
partial_product_2(39) <= temp_mult_1(39);
partial_product_2(40) <= temp_mult_1(40);
partial_product_2(41) <= temp_mult_1(41);
partial_product_2(42) <= temp_mult_1(42);
partial_product_2(43) <= temp_mult_1(43);
partial_product_2(44) <= temp_mult_1(44);
partial_product_2(45) <= temp_mult_1(45);
partial_product_2(46) <= temp_mult_1(46);
partial_product_2(47) <= temp_mult_1(47);
partial_product_2(48) <= temp_mult_1(48);
partial_product_2(49) <= temp_mult_1(49);
partial_product_2(50) <= temp_mult_1(50);
partial_product_2(51) <= temp_mult_1(51);
partial_product_2(52) <= temp_mult_1(52);
partial_product_2(53) <= temp_mult_1(53);
partial_product_2(54) <= temp_mult_1(54);
partial_product_2(55) <= temp_mult_1(55);
partial_product_2(56) <= temp_mult_1(56);
partial_product_2(57) <= temp_mult_1(57);
partial_product_2(58) <= temp_mult_1(58);
partial_product_2(59) <= temp_mult_1(59);
partial_product_2(60) <= temp_mult_1(60);
partial_product_2(61) <= temp_mult_1(61);
partial_product_2(62) <= temp_mult_1(62);
partial_product_2(63) <= temp_mult_1(63);
partial_product_2(64) <= temp_mult_1(64);
partial_product_2(65) <= temp_mult_7(65);
partial_product_2(66) <= temp_mult_7(66);
partial_product_2(67) <= temp_mult_7(67);
partial_product_2(68) <= temp_mult_7(68);
partial_product_2(69) <= temp_mult_7(69);
partial_product_2(70) <= temp_mult_7(70);
partial_product_2(71) <= temp_mult_7(71);
partial_product_2(72) <= temp_mult_7(72);
partial_product_2(73) <= temp_mult_7(73);
partial_product_2(74) <= temp_mult_7(74);
partial_product_2(75) <= temp_mult_7(75);
partial_product_2(76) <= temp_mult_7(76);
partial_product_2(77) <= temp_mult_7(77);
partial_product_2(78) <= temp_mult_7(78);
partial_product_2(79) <= temp_mult_7(79);
partial_product_2(80) <= temp_mult_7(80);
partial_product_2(81) <= temp_mult_7(81);
partial_product_2(82) <= temp_mult_7(82);
partial_product_2(83) <= temp_mult_7(83);
partial_product_2(84) <= temp_mult_7(84);
partial_product_2(85) <= temp_mult_7(85);
partial_product_2(86) <= temp_mult_7(86);
partial_product_2(87) <= temp_mult_7(87);
partial_product_2(88) <= temp_mult_7(88);
partial_product_2(89) <= temp_mult_7(89);
partial_product_2(90) <= temp_mult_7(90);
partial_product_2(91) <= temp_mult_7(91);
partial_product_2(92) <= temp_mult_7(92);
partial_product_2(93) <= temp_mult_7(93);
partial_product_2(94) <= temp_mult_7(94);
partial_product_2(95) <= temp_mult_7(95);
partial_product_2(96) <= temp_mult_7(96);
partial_product_2(97) <= temp_mult_7(97);
partial_product_2(98) <= temp_mult_7(98);
partial_product_2(99) <= temp_mult_7(99);
partial_product_2(100) <= temp_mult_7(100);
partial_product_2(101) <= temp_mult_7(101);
partial_product_2(102) <= temp_mult_7(102);
partial_product_2(103) <= temp_mult_7(103);
partial_product_2(104) <= temp_mult_7(104);
partial_product_2(105) <= temp_mult_7(105);
partial_product_2(106) <= temp_mult_13(106);
partial_product_2(107) <= temp_mult_13(107);
partial_product_2(108) <= temp_mult_13(108);
partial_product_2(109) <= temp_mult_13(109);
partial_product_2(110) <= temp_mult_13(110);
partial_product_2(111) <= temp_mult_13(111);
partial_product_2(112) <= temp_mult_13(112);
partial_product_2(113) <= temp_mult_13(113);
partial_product_2(114) <= temp_mult_13(114);
partial_product_2(115) <= temp_mult_13(115);
partial_product_2(116) <= temp_mult_13(116);
partial_product_2(117) <= temp_mult_13(117);
partial_product_2(118) <= temp_mult_13(118);
partial_product_2(119) <= temp_mult_13(119);
partial_product_2(120) <= temp_mult_13(120);
partial_product_2(121) <= temp_mult_13(121);
partial_product_2(122) <= temp_mult_13(122);
partial_product_2(123) <= temp_mult_13(123);
partial_product_2(124) <= temp_mult_13(124);
partial_product_2(125) <= temp_mult_13(125);
partial_product_2(126) <= temp_mult_13(126);
partial_product_2(127) <= temp_mult_13(127);
partial_product_2(128) <= temp_mult_13(128);
partial_product_2(129) <= temp_mult_13(129);
partial_product_2(130) <= temp_mult_13(130);
partial_product_2(131) <= temp_mult_13(131);
partial_product_2(132) <= temp_mult_13(132);
partial_product_2(133) <= temp_mult_13(133);
partial_product_2(134) <= temp_mult_13(134);
partial_product_2(135) <= temp_mult_13(135);
partial_product_2(136) <= temp_mult_13(136);
partial_product_2(137) <= temp_mult_13(137);
partial_product_2(138) <= temp_mult_13(138);
partial_product_2(139) <= temp_mult_13(139);
partial_product_2(140) <= temp_mult_13(140);
partial_product_2(141) <= temp_mult_13(141);
partial_product_2(142) <= temp_mult_13(142);
partial_product_2(143) <= temp_mult_13(143);
partial_product_2(144) <= temp_mult_13(144);
partial_product_2(145) <= temp_mult_13(145);
partial_product_2(146) <= temp_mult_13(146);
partial_product_2(147) <= temp_mult_19(147);
partial_product_2(148) <= temp_mult_19(148);
partial_product_2(149) <= temp_mult_19(149);
partial_product_2(150) <= temp_mult_19(150);
partial_product_2(151) <= temp_mult_19(151);
partial_product_2(152) <= temp_mult_19(152);
partial_product_2(153) <= temp_mult_19(153);
partial_product_2(154) <= temp_mult_19(154);
partial_product_2(155) <= temp_mult_19(155);
partial_product_2(156) <= temp_mult_19(156);
partial_product_2(157) <= temp_mult_19(157);
partial_product_2(158) <= temp_mult_19(158);
partial_product_2(159) <= temp_mult_19(159);
partial_product_2(160) <= temp_mult_19(160);
partial_product_2(161) <= temp_mult_19(161);
partial_product_2(162) <= temp_mult_19(162);
partial_product_2(163) <= temp_mult_19(163);
partial_product_2(164) <= temp_mult_19(164);
partial_product_2(165) <= temp_mult_19(165);
partial_product_2(166) <= temp_mult_19(166);
partial_product_2(167) <= temp_mult_19(167);
partial_product_2(168) <= temp_mult_19(168);
partial_product_2(169) <= temp_mult_19(169);
partial_product_2(170) <= temp_mult_19(170);
partial_product_2(171) <= temp_mult_19(171);
partial_product_2(172) <= temp_mult_19(172);
partial_product_2(173) <= temp_mult_19(173);
partial_product_2(174) <= temp_mult_19(174);
partial_product_2(175) <= temp_mult_19(175);
partial_product_2(176) <= temp_mult_19(176);
partial_product_2(177) <= temp_mult_19(177);
partial_product_2(178) <= temp_mult_19(178);
partial_product_2(179) <= temp_mult_19(179);
partial_product_2(180) <= temp_mult_19(180);
partial_product_2(181) <= temp_mult_19(181);
partial_product_2(182) <= temp_mult_19(182);
partial_product_2(183) <= temp_mult_19(183);
partial_product_2(184) <= temp_mult_19(184);
partial_product_2(185) <= temp_mult_19(185);
partial_product_2(186) <= temp_mult_19(186);
partial_product_2(187) <= temp_mult_19(187);
partial_product_2(188) <= temp_mult_44(188);
partial_product_2(189) <= temp_mult_44(189);
partial_product_2(190) <= temp_mult_44(190);
partial_product_2(191) <= temp_mult_44(191);
partial_product_2(192) <= temp_mult_44(192);
partial_product_2(193) <= temp_mult_44(193);
partial_product_2(194) <= temp_mult_44(194);
partial_product_2(195) <= temp_mult_44(195);
partial_product_2(196) <= temp_mult_44(196);
partial_product_2(197) <= temp_mult_44(197);
partial_product_2(198) <= temp_mult_44(198);
partial_product_2(199) <= temp_mult_44(199);
partial_product_2(200) <= temp_mult_44(200);
partial_product_2(201) <= temp_mult_44(201);
partial_product_2(202) <= temp_mult_44(202);
partial_product_2(203) <= temp_mult_44(203);
partial_product_2(204) <= temp_mult_44(204);
partial_product_2(205) <= temp_mult_44(205);
partial_product_2(206) <= temp_mult_44(206);
partial_product_2(207) <= temp_mult_44(207);
partial_product_2(208) <= temp_mult_44(208);
partial_product_2(209) <= temp_mult_44(209);
partial_product_2(210) <= temp_mult_44(210);
partial_product_2(211) <= temp_mult_44(211);
partial_product_2(212) <= temp_mult_44(212);
partial_product_2(213) <= temp_mult_44(213);
partial_product_2(214) <= temp_mult_44(214);
partial_product_2(215) <= temp_mult_44(215);
partial_product_2(216) <= temp_mult_44(216);
partial_product_2(217) <= temp_mult_44(217);
partial_product_2(218) <= temp_mult_44(218);
partial_product_2(219) <= temp_mult_44(219);
partial_product_2(220) <= temp_mult_44(220);
partial_product_2(221) <= temp_mult_44(221);
partial_product_2(222) <= temp_mult_44(222);
partial_product_2(223) <= temp_mult_44(223);
partial_product_2(224) <= temp_mult_44(224);
partial_product_2(225) <= temp_mult_44(225);
partial_product_2(226) <= temp_mult_44(226);
partial_product_2(227) <= temp_mult_44(227);
partial_product_2(228) <= temp_mult_44(228);
partial_product_2(229) <= temp_mult_53(229);
partial_product_2(230) <= temp_mult_53(230);
partial_product_2(231) <= temp_mult_53(231);
partial_product_2(232) <= temp_mult_53(232);
partial_product_2(233) <= temp_mult_53(233);
partial_product_2(234) <= temp_mult_53(234);
partial_product_2(235) <= temp_mult_53(235);
partial_product_2(236) <= temp_mult_53(236);
partial_product_2(237) <= temp_mult_53(237);
partial_product_2(238) <= temp_mult_53(238);
partial_product_2(239) <= temp_mult_53(239);
partial_product_2(240) <= temp_mult_53(240);
partial_product_2(241) <= temp_mult_53(241);
partial_product_2(242) <= temp_mult_53(242);
partial_product_2(243) <= temp_mult_53(243);
partial_product_2(244) <= temp_mult_53(244);
partial_product_2(245) <= temp_mult_53(245);
partial_product_2(246) <= temp_mult_53(246);
partial_product_2(247) <= temp_mult_53(247);
partial_product_2(248) <= temp_mult_53(248);
partial_product_2(249) <= temp_mult_53(249);
partial_product_2(250) <= temp_mult_53(250);
partial_product_2(251) <= temp_mult_53(251);
partial_product_2(252) <= temp_mult_53(252);
partial_product_2(253) <= temp_mult_53(253);
partial_product_2(254) <= temp_mult_53(254);
partial_product_2(255) <= temp_mult_53(255);
partial_product_2(256) <= temp_mult_53(256);
partial_product_2(257) <= temp_mult_53(257);
partial_product_2(258) <= temp_mult_53(258);
partial_product_2(259) <= temp_mult_53(259);
partial_product_2(260) <= temp_mult_53(260);
partial_product_2(261) <= temp_mult_53(261);
partial_product_2(262) <= temp_mult_53(262);
partial_product_2(263) <= temp_mult_53(263);
partial_product_2(264) <= temp_mult_53(264);
partial_product_2(265) <= temp_mult_53(265);
partial_product_2(266) <= temp_mult_53(266);
partial_product_2(267) <= temp_mult_53(267);
partial_product_2(268) <= temp_mult_53(268);
partial_product_2(269) <= temp_mult_53(269);
partial_product_2(270) <= temp_mult_62(270);
partial_product_2(271) <= temp_mult_62(271);
partial_product_2(272) <= temp_mult_62(272);
partial_product_2(273) <= temp_mult_62(273);
partial_product_2(274) <= temp_mult_62(274);
partial_product_2(275) <= temp_mult_62(275);
partial_product_2(276) <= temp_mult_62(276);
partial_product_2(277) <= temp_mult_62(277);
partial_product_2(278) <= temp_mult_62(278);
partial_product_2(279) <= temp_mult_62(279);
partial_product_2(280) <= temp_mult_62(280);
partial_product_2(281) <= temp_mult_62(281);
partial_product_2(282) <= temp_mult_62(282);
partial_product_2(283) <= temp_mult_62(283);
partial_product_2(284) <= temp_mult_62(284);
partial_product_2(285) <= temp_mult_62(285);
partial_product_2(286) <= temp_mult_62(286);
partial_product_2(287) <= temp_mult_62(287);
partial_product_2(288) <= temp_mult_62(288);
partial_product_2(289) <= temp_mult_62(289);
partial_product_2(290) <= temp_mult_62(290);
partial_product_2(291) <= temp_mult_62(291);
partial_product_2(292) <= temp_mult_62(292);
partial_product_2(293) <= temp_mult_62(293);
partial_product_2(294) <= temp_mult_62(294);
partial_product_2(295) <= temp_mult_62(295);
partial_product_2(296) <= temp_mult_62(296);
partial_product_2(297) <= temp_mult_62(297);
partial_product_2(298) <= temp_mult_62(298);
partial_product_2(299) <= temp_mult_62(299);
partial_product_2(300) <= temp_mult_62(300);
partial_product_2(301) <= temp_mult_62(301);
partial_product_2(302) <= temp_mult_62(302);
partial_product_2(303) <= temp_mult_62(303);
partial_product_2(304) <= temp_mult_62(304);
partial_product_2(305) <= temp_mult_62(305);
partial_product_2(306) <= temp_mult_62(306);
partial_product_2(307) <= temp_mult_62(307);
partial_product_2(308) <= temp_mult_62(308);
partial_product_2(309) <= temp_mult_62(309);
partial_product_2(310) <= temp_mult_62(310);
partial_product_2(311) <= temp_mult_71(311);
partial_product_2(312) <= temp_mult_71(312);
partial_product_2(313) <= temp_mult_71(313);
partial_product_2(314) <= temp_mult_71(314);
partial_product_2(315) <= temp_mult_71(315);
partial_product_2(316) <= temp_mult_71(316);
partial_product_2(317) <= temp_mult_71(317);
partial_product_2(318) <= temp_mult_71(318);
partial_product_2(319) <= temp_mult_71(319);
partial_product_2(320) <= temp_mult_71(320);
partial_product_2(321) <= temp_mult_71(321);
partial_product_2(322) <= temp_mult_71(322);
partial_product_2(323) <= temp_mult_71(323);
partial_product_2(324) <= temp_mult_71(324);
partial_product_2(325) <= temp_mult_71(325);
partial_product_2(326) <= temp_mult_71(326);
partial_product_2(327) <= temp_mult_71(327);
partial_product_2(328) <= temp_mult_71(328);
partial_product_2(329) <= temp_mult_71(329);
partial_product_2(330) <= temp_mult_71(330);
partial_product_2(331) <= temp_mult_71(331);
partial_product_2(332) <= temp_mult_71(332);
partial_product_2(333) <= temp_mult_71(333);
partial_product_2(334) <= temp_mult_71(334);
partial_product_2(335) <= temp_mult_71(335);
partial_product_2(336) <= temp_mult_71(336);
partial_product_2(337) <= temp_mult_71(337);
partial_product_2(338) <= temp_mult_71(338);
partial_product_2(339) <= temp_mult_71(339);
partial_product_2(340) <= temp_mult_71(340);
partial_product_2(341) <= temp_mult_71(341);
partial_product_2(342) <= temp_mult_71(342);
partial_product_2(343) <= temp_mult_71(343);
partial_product_2(344) <= temp_mult_71(344);
partial_product_2(345) <= temp_mult_71(345);
partial_product_2(346) <= temp_mult_71(346);
partial_product_2(347) <= temp_mult_71(347);
partial_product_2(348) <= temp_mult_71(348);
partial_product_2(349) <= temp_mult_71(349);
partial_product_2(350) <= temp_mult_71(350);
partial_product_2(351) <= temp_mult_71(351);
partial_product_2(352) <= temp_mult_124(352);
partial_product_2(353) <= temp_mult_124(353);
partial_product_2(354) <= temp_mult_124(354);
partial_product_2(355) <= temp_mult_124(355);
partial_product_2(356) <= temp_mult_124(356);
partial_product_2(357) <= temp_mult_124(357);
partial_product_2(358) <= temp_mult_124(358);
partial_product_2(359) <= temp_mult_124(359);
partial_product_2(360) <= temp_mult_124(360);
partial_product_2(361) <= temp_mult_124(361);
partial_product_2(362) <= temp_mult_124(362);
partial_product_2(363) <= temp_mult_124(363);
partial_product_2(364) <= temp_mult_124(364);
partial_product_2(365) <= temp_mult_124(365);
partial_product_2(366) <= temp_mult_124(366);
partial_product_2(367) <= temp_mult_124(367);
partial_product_2(368) <= temp_mult_124(368);
partial_product_2(369) <= temp_mult_124(369);
partial_product_2(370) <= temp_mult_124(370);
partial_product_2(371) <= temp_mult_124(371);
partial_product_2(372) <= temp_mult_124(372);
partial_product_2(373) <= temp_mult_124(373);
partial_product_2(374) <= temp_mult_124(374);
partial_product_2(375) <= temp_mult_124(375);
partial_product_2(376) <= temp_mult_124(376);
partial_product_2(377) <= temp_mult_124(377);
partial_product_2(378) <= temp_mult_124(378);
partial_product_2(379) <= temp_mult_124(379);
partial_product_2(380) <= temp_mult_124(380);
partial_product_2(381) <= temp_mult_124(381);
partial_product_2(382) <= temp_mult_124(382);
partial_product_2(383) <= temp_mult_124(383);
partial_product_2(384) <= temp_mult_124(384);
partial_product_2(385) <= temp_mult_124(385);
partial_product_2(386) <= temp_mult_124(386);
partial_product_2(387) <= temp_mult_124(387);
partial_product_2(388) <= temp_mult_124(388);
partial_product_2(389) <= temp_mult_124(389);
partial_product_2(390) <= temp_mult_124(390);
partial_product_2(391) <= temp_mult_124(391);
partial_product_2(392) <= temp_mult_124(392);
partial_product_2(393) <= '0';
partial_product_2(394) <= '0';
partial_product_2(395) <= '0';
partial_product_2(396) <= temp_mult_143(396);
partial_product_2(397) <= temp_mult_143(397);
partial_product_2(398) <= temp_mult_143(398);
partial_product_2(399) <= temp_mult_143(399);
partial_product_2(400) <= temp_mult_143(400);
partial_product_2(401) <= temp_mult_143(401);
partial_product_2(402) <= temp_mult_143(402);
partial_product_2(403) <= temp_mult_143(403);
partial_product_2(404) <= temp_mult_143(404);
partial_product_2(405) <= temp_mult_143(405);
partial_product_2(406) <= temp_mult_143(406);
partial_product_2(407) <= temp_mult_143(407);
partial_product_2(408) <= temp_mult_143(408);
partial_product_2(409) <= temp_mult_143(409);
partial_product_2(410) <= temp_mult_143(410);
partial_product_2(411) <= temp_mult_143(411);
partial_product_2(412) <= temp_mult_143(412);
partial_product_2(413) <= temp_mult_143(413);
partial_product_2(414) <= temp_mult_143(414);
partial_product_2(415) <= temp_mult_143(415);
partial_product_2(416) <= temp_mult_143(416);
partial_product_2(417) <= temp_mult_143(417);
partial_product_2(418) <= temp_mult_143(418);
partial_product_2(419) <= temp_mult_143(419);
partial_product_2(420) <= temp_mult_143(420);
partial_product_2(421) <= temp_mult_143(421);
partial_product_2(422) <= temp_mult_143(422);
partial_product_2(423) <= temp_mult_143(423);
partial_product_2(424) <= temp_mult_143(424);
partial_product_2(425) <= temp_mult_143(425);
partial_product_2(426) <= temp_mult_143(426);
partial_product_2(427) <= temp_mult_143(427);
partial_product_2(428) <= temp_mult_143(428);
partial_product_2(429) <= temp_mult_143(429);
partial_product_2(430) <= temp_mult_143(430);
partial_product_2(431) <= temp_mult_143(431);
partial_product_2(432) <= temp_mult_143(432);
partial_product_2(433) <= temp_mult_143(433);
partial_product_2(434) <= temp_mult_143(434);
partial_product_2(435) <= temp_mult_143(435);
partial_product_2(436) <= temp_mult_143(436);
partial_product_2(437) <= temp_mult_149(437);
partial_product_2(438) <= temp_mult_149(438);
partial_product_2(439) <= temp_mult_149(439);
partial_product_2(440) <= temp_mult_149(440);
partial_product_2(441) <= temp_mult_149(441);
partial_product_2(442) <= temp_mult_149(442);
partial_product_2(443) <= temp_mult_149(443);
partial_product_2(444) <= temp_mult_149(444);
partial_product_2(445) <= temp_mult_149(445);
partial_product_2(446) <= temp_mult_149(446);
partial_product_2(447) <= temp_mult_149(447);
partial_product_2(448) <= temp_mult_149(448);
partial_product_2(449) <= temp_mult_149(449);
partial_product_2(450) <= temp_mult_149(450);
partial_product_2(451) <= temp_mult_149(451);
partial_product_2(452) <= temp_mult_149(452);
partial_product_2(453) <= temp_mult_149(453);
partial_product_2(454) <= temp_mult_149(454);
partial_product_2(455) <= temp_mult_149(455);
partial_product_2(456) <= temp_mult_149(456);
partial_product_2(457) <= temp_mult_149(457);
partial_product_2(458) <= temp_mult_149(458);
partial_product_2(459) <= temp_mult_149(459);
partial_product_2(460) <= temp_mult_149(460);
partial_product_2(461) <= temp_mult_149(461);
partial_product_2(462) <= temp_mult_149(462);
partial_product_2(463) <= temp_mult_149(463);
partial_product_2(464) <= temp_mult_149(464);
partial_product_2(465) <= temp_mult_149(465);
partial_product_2(466) <= temp_mult_149(466);
partial_product_2(467) <= temp_mult_149(467);
partial_product_2(468) <= temp_mult_149(468);
partial_product_2(469) <= temp_mult_149(469);
partial_product_2(470) <= temp_mult_149(470);
partial_product_2(471) <= temp_mult_149(471);
partial_product_2(472) <= temp_mult_149(472);
partial_product_2(473) <= temp_mult_149(473);
partial_product_2(474) <= temp_mult_149(474);
partial_product_2(475) <= temp_mult_149(475);
partial_product_2(476) <= temp_mult_149(476);
partial_product_2(477) <= temp_mult_149(477);
partial_product_2(478) <= '0';
partial_product_2(479) <= '0';
partial_product_2(480) <= '0';
partial_product_2(481) <= '0';
partial_product_2(482) <= '0';
partial_product_2(483) <= '0';
partial_product_2(484) <= '0';
partial_product_2(485) <= '0';
partial_product_2(486) <= '0';
partial_product_2(487) <= '0';
partial_product_2(488) <= '0';
partial_product_2(489) <= '0';
partial_product_2(490) <= '0';
partial_product_2(491) <= '0';
partial_product_2(492) <= '0';
partial_product_2(493) <= '0';
partial_product_2(494) <= '0';
partial_product_2(495) <= '0';
partial_product_2(496) <= '0';
partial_product_2(497) <= '0';
partial_product_2(498) <= '0';
partial_product_2(499) <= '0';
partial_product_2(500) <= '0';
partial_product_2(501) <= '0';
partial_product_2(502) <= '0';
partial_product_2(503) <= '0';
partial_product_2(504) <= '0';
partial_product_2(505) <= '0';
partial_product_2(506) <= '0';
partial_product_2(507) <= '0';
partial_product_2(508) <= '0';
partial_product_2(509) <= '0';
partial_product_2(510) <= '0';
partial_product_2(511) <= '0';
partial_product_2(512) <= '0';
partial_product_3(0) <= '0';
partial_product_3(1) <= '0';
partial_product_3(2) <= '0';
partial_product_3(3) <= '0';
partial_product_3(4) <= '0';
partial_product_3(5) <= '0';
partial_product_3(6) <= '0';
partial_product_3(7) <= '0';
partial_product_3(8) <= '0';
partial_product_3(9) <= '0';
partial_product_3(10) <= '0';
partial_product_3(11) <= '0';
partial_product_3(12) <= '0';
partial_product_3(13) <= '0';
partial_product_3(14) <= '0';
partial_product_3(15) <= '0';
partial_product_3(16) <= '0';
partial_product_3(17) <= '0';
partial_product_3(18) <= '0';
partial_product_3(19) <= '0';
partial_product_3(20) <= '0';
partial_product_3(21) <= '0';
partial_product_3(22) <= '0';
partial_product_3(23) <= '0';
partial_product_3(24) <= '0';
partial_product_3(25) <= '0';
partial_product_3(26) <= '0';
partial_product_3(27) <= '0';
partial_product_3(28) <= '0';
partial_product_3(29) <= '0';
partial_product_3(30) <= '0';
partial_product_3(31) <= '0';
partial_product_3(32) <= '0';
partial_product_3(33) <= '0';
partial_product_3(34) <= temp_mult_10(34);
partial_product_3(35) <= temp_mult_10(35);
partial_product_3(36) <= temp_mult_10(36);
partial_product_3(37) <= temp_mult_10(37);
partial_product_3(38) <= temp_mult_10(38);
partial_product_3(39) <= temp_mult_10(39);
partial_product_3(40) <= temp_mult_10(40);
partial_product_3(41) <= temp_mult_10(41);
partial_product_3(42) <= temp_mult_10(42);
partial_product_3(43) <= temp_mult_10(43);
partial_product_3(44) <= temp_mult_10(44);
partial_product_3(45) <= temp_mult_10(45);
partial_product_3(46) <= temp_mult_10(46);
partial_product_3(47) <= temp_mult_10(47);
partial_product_3(48) <= temp_mult_10(48);
partial_product_3(49) <= temp_mult_10(49);
partial_product_3(50) <= temp_mult_10(50);
partial_product_3(51) <= temp_mult_10(51);
partial_product_3(52) <= temp_mult_10(52);
partial_product_3(53) <= temp_mult_10(53);
partial_product_3(54) <= temp_mult_10(54);
partial_product_3(55) <= temp_mult_10(55);
partial_product_3(56) <= temp_mult_10(56);
partial_product_3(57) <= temp_mult_10(57);
partial_product_3(58) <= temp_mult_10(58);
partial_product_3(59) <= temp_mult_10(59);
partial_product_3(60) <= temp_mult_10(60);
partial_product_3(61) <= temp_mult_10(61);
partial_product_3(62) <= temp_mult_10(62);
partial_product_3(63) <= temp_mult_10(63);
partial_product_3(64) <= temp_mult_10(64);
partial_product_3(65) <= temp_mult_10(65);
partial_product_3(66) <= temp_mult_10(66);
partial_product_3(67) <= temp_mult_10(67);
partial_product_3(68) <= temp_mult_10(68);
partial_product_3(69) <= temp_mult_10(69);
partial_product_3(70) <= temp_mult_10(70);
partial_product_3(71) <= temp_mult_10(71);
partial_product_3(72) <= temp_mult_10(72);
partial_product_3(73) <= temp_mult_10(73);
partial_product_3(74) <= temp_mult_10(74);
partial_product_3(75) <= temp_mult_16(75);
partial_product_3(76) <= temp_mult_16(76);
partial_product_3(77) <= temp_mult_16(77);
partial_product_3(78) <= temp_mult_16(78);
partial_product_3(79) <= temp_mult_16(79);
partial_product_3(80) <= temp_mult_16(80);
partial_product_3(81) <= temp_mult_16(81);
partial_product_3(82) <= temp_mult_16(82);
partial_product_3(83) <= temp_mult_16(83);
partial_product_3(84) <= temp_mult_16(84);
partial_product_3(85) <= temp_mult_16(85);
partial_product_3(86) <= temp_mult_16(86);
partial_product_3(87) <= temp_mult_16(87);
partial_product_3(88) <= temp_mult_16(88);
partial_product_3(89) <= temp_mult_16(89);
partial_product_3(90) <= temp_mult_16(90);
partial_product_3(91) <= temp_mult_16(91);
partial_product_3(92) <= temp_mult_16(92);
partial_product_3(93) <= temp_mult_16(93);
partial_product_3(94) <= temp_mult_16(94);
partial_product_3(95) <= temp_mult_16(95);
partial_product_3(96) <= temp_mult_16(96);
partial_product_3(97) <= temp_mult_16(97);
partial_product_3(98) <= temp_mult_16(98);
partial_product_3(99) <= temp_mult_16(99);
partial_product_3(100) <= temp_mult_16(100);
partial_product_3(101) <= temp_mult_16(101);
partial_product_3(102) <= temp_mult_16(102);
partial_product_3(103) <= temp_mult_16(103);
partial_product_3(104) <= temp_mult_16(104);
partial_product_3(105) <= temp_mult_16(105);
partial_product_3(106) <= temp_mult_16(106);
partial_product_3(107) <= temp_mult_16(107);
partial_product_3(108) <= temp_mult_16(108);
partial_product_3(109) <= temp_mult_16(109);
partial_product_3(110) <= temp_mult_16(110);
partial_product_3(111) <= temp_mult_16(111);
partial_product_3(112) <= temp_mult_16(112);
partial_product_3(113) <= temp_mult_16(113);
partial_product_3(114) <= temp_mult_16(114);
partial_product_3(115) <= temp_mult_16(115);
partial_product_3(116) <= temp_mult_22(116);
partial_product_3(117) <= temp_mult_22(117);
partial_product_3(118) <= temp_mult_22(118);
partial_product_3(119) <= temp_mult_22(119);
partial_product_3(120) <= temp_mult_22(120);
partial_product_3(121) <= temp_mult_22(121);
partial_product_3(122) <= temp_mult_22(122);
partial_product_3(123) <= temp_mult_22(123);
partial_product_3(124) <= temp_mult_22(124);
partial_product_3(125) <= temp_mult_22(125);
partial_product_3(126) <= temp_mult_22(126);
partial_product_3(127) <= temp_mult_22(127);
partial_product_3(128) <= temp_mult_22(128);
partial_product_3(129) <= temp_mult_22(129);
partial_product_3(130) <= temp_mult_22(130);
partial_product_3(131) <= temp_mult_22(131);
partial_product_3(132) <= temp_mult_22(132);
partial_product_3(133) <= temp_mult_22(133);
partial_product_3(134) <= temp_mult_22(134);
partial_product_3(135) <= temp_mult_22(135);
partial_product_3(136) <= temp_mult_22(136);
partial_product_3(137) <= temp_mult_22(137);
partial_product_3(138) <= temp_mult_22(138);
partial_product_3(139) <= temp_mult_22(139);
partial_product_3(140) <= temp_mult_22(140);
partial_product_3(141) <= temp_mult_22(141);
partial_product_3(142) <= temp_mult_22(142);
partial_product_3(143) <= temp_mult_22(143);
partial_product_3(144) <= temp_mult_22(144);
partial_product_3(145) <= temp_mult_22(145);
partial_product_3(146) <= temp_mult_22(146);
partial_product_3(147) <= temp_mult_22(147);
partial_product_3(148) <= temp_mult_22(148);
partial_product_3(149) <= temp_mult_22(149);
partial_product_3(150) <= temp_mult_22(150);
partial_product_3(151) <= temp_mult_22(151);
partial_product_3(152) <= temp_mult_22(152);
partial_product_3(153) <= temp_mult_22(153);
partial_product_3(154) <= temp_mult_22(154);
partial_product_3(155) <= temp_mult_22(155);
partial_product_3(156) <= temp_mult_22(156);
partial_product_3(157) <= temp_mult_28(157);
partial_product_3(158) <= temp_mult_28(158);
partial_product_3(159) <= temp_mult_28(159);
partial_product_3(160) <= temp_mult_28(160);
partial_product_3(161) <= temp_mult_28(161);
partial_product_3(162) <= temp_mult_28(162);
partial_product_3(163) <= temp_mult_28(163);
partial_product_3(164) <= temp_mult_28(164);
partial_product_3(165) <= temp_mult_28(165);
partial_product_3(166) <= temp_mult_28(166);
partial_product_3(167) <= temp_mult_28(167);
partial_product_3(168) <= temp_mult_28(168);
partial_product_3(169) <= temp_mult_28(169);
partial_product_3(170) <= temp_mult_28(170);
partial_product_3(171) <= temp_mult_28(171);
partial_product_3(172) <= temp_mult_28(172);
partial_product_3(173) <= temp_mult_28(173);
partial_product_3(174) <= temp_mult_28(174);
partial_product_3(175) <= temp_mult_28(175);
partial_product_3(176) <= temp_mult_28(176);
partial_product_3(177) <= temp_mult_28(177);
partial_product_3(178) <= temp_mult_28(178);
partial_product_3(179) <= temp_mult_28(179);
partial_product_3(180) <= temp_mult_28(180);
partial_product_3(181) <= temp_mult_28(181);
partial_product_3(182) <= temp_mult_28(182);
partial_product_3(183) <= temp_mult_28(183);
partial_product_3(184) <= temp_mult_28(184);
partial_product_3(185) <= temp_mult_28(185);
partial_product_3(186) <= temp_mult_28(186);
partial_product_3(187) <= temp_mult_28(187);
partial_product_3(188) <= temp_mult_28(188);
partial_product_3(189) <= temp_mult_28(189);
partial_product_3(190) <= temp_mult_28(190);
partial_product_3(191) <= temp_mult_28(191);
partial_product_3(192) <= temp_mult_28(192);
partial_product_3(193) <= temp_mult_28(193);
partial_product_3(194) <= temp_mult_28(194);
partial_product_3(195) <= temp_mult_28(195);
partial_product_3(196) <= temp_mult_28(196);
partial_product_3(197) <= temp_mult_28(197);
partial_product_3(198) <= temp_mult_34(198);
partial_product_3(199) <= temp_mult_34(199);
partial_product_3(200) <= temp_mult_34(200);
partial_product_3(201) <= temp_mult_34(201);
partial_product_3(202) <= temp_mult_34(202);
partial_product_3(203) <= temp_mult_34(203);
partial_product_3(204) <= temp_mult_34(204);
partial_product_3(205) <= temp_mult_34(205);
partial_product_3(206) <= temp_mult_34(206);
partial_product_3(207) <= temp_mult_34(207);
partial_product_3(208) <= temp_mult_34(208);
partial_product_3(209) <= temp_mult_34(209);
partial_product_3(210) <= temp_mult_34(210);
partial_product_3(211) <= temp_mult_34(211);
partial_product_3(212) <= temp_mult_34(212);
partial_product_3(213) <= temp_mult_34(213);
partial_product_3(214) <= temp_mult_34(214);
partial_product_3(215) <= temp_mult_34(215);
partial_product_3(216) <= temp_mult_34(216);
partial_product_3(217) <= temp_mult_34(217);
partial_product_3(218) <= temp_mult_34(218);
partial_product_3(219) <= temp_mult_34(219);
partial_product_3(220) <= temp_mult_34(220);
partial_product_3(221) <= temp_mult_34(221);
partial_product_3(222) <= temp_mult_34(222);
partial_product_3(223) <= temp_mult_34(223);
partial_product_3(224) <= temp_mult_34(224);
partial_product_3(225) <= temp_mult_34(225);
partial_product_3(226) <= temp_mult_34(226);
partial_product_3(227) <= temp_mult_34(227);
partial_product_3(228) <= temp_mult_34(228);
partial_product_3(229) <= temp_mult_34(229);
partial_product_3(230) <= temp_mult_34(230);
partial_product_3(231) <= temp_mult_34(231);
partial_product_3(232) <= temp_mult_34(232);
partial_product_3(233) <= temp_mult_34(233);
partial_product_3(234) <= temp_mult_34(234);
partial_product_3(235) <= temp_mult_34(235);
partial_product_3(236) <= temp_mult_34(236);
partial_product_3(237) <= temp_mult_34(237);
partial_product_3(238) <= temp_mult_34(238);
partial_product_3(239) <= temp_mult_47(239);
partial_product_3(240) <= temp_mult_47(240);
partial_product_3(241) <= temp_mult_47(241);
partial_product_3(242) <= temp_mult_47(242);
partial_product_3(243) <= temp_mult_47(243);
partial_product_3(244) <= temp_mult_47(244);
partial_product_3(245) <= temp_mult_47(245);
partial_product_3(246) <= temp_mult_47(246);
partial_product_3(247) <= temp_mult_47(247);
partial_product_3(248) <= temp_mult_47(248);
partial_product_3(249) <= temp_mult_47(249);
partial_product_3(250) <= temp_mult_47(250);
partial_product_3(251) <= temp_mult_47(251);
partial_product_3(252) <= temp_mult_47(252);
partial_product_3(253) <= temp_mult_47(253);
partial_product_3(254) <= temp_mult_47(254);
partial_product_3(255) <= temp_mult_47(255);
partial_product_3(256) <= temp_mult_47(256);
partial_product_3(257) <= temp_mult_47(257);
partial_product_3(258) <= temp_mult_47(258);
partial_product_3(259) <= temp_mult_47(259);
partial_product_3(260) <= temp_mult_47(260);
partial_product_3(261) <= temp_mult_47(261);
partial_product_3(262) <= temp_mult_47(262);
partial_product_3(263) <= temp_mult_47(263);
partial_product_3(264) <= temp_mult_47(264);
partial_product_3(265) <= temp_mult_47(265);
partial_product_3(266) <= temp_mult_47(266);
partial_product_3(267) <= temp_mult_47(267);
partial_product_3(268) <= temp_mult_47(268);
partial_product_3(269) <= temp_mult_47(269);
partial_product_3(270) <= temp_mult_47(270);
partial_product_3(271) <= temp_mult_47(271);
partial_product_3(272) <= temp_mult_47(272);
partial_product_3(273) <= temp_mult_47(273);
partial_product_3(274) <= temp_mult_47(274);
partial_product_3(275) <= temp_mult_47(275);
partial_product_3(276) <= temp_mult_47(276);
partial_product_3(277) <= temp_mult_47(277);
partial_product_3(278) <= temp_mult_47(278);
partial_product_3(279) <= temp_mult_47(279);
partial_product_3(280) <= temp_mult_121(280);
partial_product_3(281) <= temp_mult_121(281);
partial_product_3(282) <= temp_mult_121(282);
partial_product_3(283) <= temp_mult_121(283);
partial_product_3(284) <= temp_mult_121(284);
partial_product_3(285) <= temp_mult_121(285);
partial_product_3(286) <= temp_mult_121(286);
partial_product_3(287) <= temp_mult_121(287);
partial_product_3(288) <= temp_mult_121(288);
partial_product_3(289) <= temp_mult_121(289);
partial_product_3(290) <= temp_mult_121(290);
partial_product_3(291) <= temp_mult_121(291);
partial_product_3(292) <= temp_mult_121(292);
partial_product_3(293) <= temp_mult_121(293);
partial_product_3(294) <= temp_mult_121(294);
partial_product_3(295) <= temp_mult_121(295);
partial_product_3(296) <= temp_mult_121(296);
partial_product_3(297) <= temp_mult_121(297);
partial_product_3(298) <= temp_mult_121(298);
partial_product_3(299) <= temp_mult_121(299);
partial_product_3(300) <= temp_mult_121(300);
partial_product_3(301) <= temp_mult_121(301);
partial_product_3(302) <= temp_mult_121(302);
partial_product_3(303) <= temp_mult_121(303);
partial_product_3(304) <= temp_mult_121(304);
partial_product_3(305) <= temp_mult_121(305);
partial_product_3(306) <= temp_mult_121(306);
partial_product_3(307) <= temp_mult_121(307);
partial_product_3(308) <= temp_mult_121(308);
partial_product_3(309) <= temp_mult_121(309);
partial_product_3(310) <= temp_mult_121(310);
partial_product_3(311) <= temp_mult_121(311);
partial_product_3(312) <= temp_mult_121(312);
partial_product_3(313) <= temp_mult_121(313);
partial_product_3(314) <= temp_mult_121(314);
partial_product_3(315) <= temp_mult_121(315);
partial_product_3(316) <= temp_mult_121(316);
partial_product_3(317) <= temp_mult_121(317);
partial_product_3(318) <= temp_mult_121(318);
partial_product_3(319) <= temp_mult_121(319);
partial_product_3(320) <= temp_mult_121(320);
partial_product_3(321) <= temp_mult_127(321);
partial_product_3(322) <= temp_mult_127(322);
partial_product_3(323) <= temp_mult_127(323);
partial_product_3(324) <= temp_mult_127(324);
partial_product_3(325) <= temp_mult_127(325);
partial_product_3(326) <= temp_mult_127(326);
partial_product_3(327) <= temp_mult_127(327);
partial_product_3(328) <= temp_mult_127(328);
partial_product_3(329) <= temp_mult_127(329);
partial_product_3(330) <= temp_mult_127(330);
partial_product_3(331) <= temp_mult_127(331);
partial_product_3(332) <= temp_mult_127(332);
partial_product_3(333) <= temp_mult_127(333);
partial_product_3(334) <= temp_mult_127(334);
partial_product_3(335) <= temp_mult_127(335);
partial_product_3(336) <= temp_mult_127(336);
partial_product_3(337) <= temp_mult_127(337);
partial_product_3(338) <= temp_mult_127(338);
partial_product_3(339) <= temp_mult_127(339);
partial_product_3(340) <= temp_mult_127(340);
partial_product_3(341) <= temp_mult_127(341);
partial_product_3(342) <= temp_mult_127(342);
partial_product_3(343) <= temp_mult_127(343);
partial_product_3(344) <= temp_mult_127(344);
partial_product_3(345) <= temp_mult_127(345);
partial_product_3(346) <= temp_mult_127(346);
partial_product_3(347) <= temp_mult_127(347);
partial_product_3(348) <= temp_mult_127(348);
partial_product_3(349) <= temp_mult_127(349);
partial_product_3(350) <= temp_mult_127(350);
partial_product_3(351) <= temp_mult_127(351);
partial_product_3(352) <= temp_mult_127(352);
partial_product_3(353) <= temp_mult_127(353);
partial_product_3(354) <= temp_mult_127(354);
partial_product_3(355) <= temp_mult_127(355);
partial_product_3(356) <= temp_mult_127(356);
partial_product_3(357) <= temp_mult_127(357);
partial_product_3(358) <= temp_mult_127(358);
partial_product_3(359) <= temp_mult_127(359);
partial_product_3(360) <= temp_mult_127(360);
partial_product_3(361) <= temp_mult_127(361);
partial_product_3(362) <= temp_mult_133(362);
partial_product_3(363) <= temp_mult_133(363);
partial_product_3(364) <= temp_mult_133(364);
partial_product_3(365) <= temp_mult_133(365);
partial_product_3(366) <= temp_mult_133(366);
partial_product_3(367) <= temp_mult_133(367);
partial_product_3(368) <= temp_mult_133(368);
partial_product_3(369) <= temp_mult_133(369);
partial_product_3(370) <= temp_mult_133(370);
partial_product_3(371) <= temp_mult_133(371);
partial_product_3(372) <= temp_mult_133(372);
partial_product_3(373) <= temp_mult_133(373);
partial_product_3(374) <= temp_mult_133(374);
partial_product_3(375) <= temp_mult_133(375);
partial_product_3(376) <= temp_mult_133(376);
partial_product_3(377) <= temp_mult_133(377);
partial_product_3(378) <= temp_mult_133(378);
partial_product_3(379) <= temp_mult_133(379);
partial_product_3(380) <= temp_mult_133(380);
partial_product_3(381) <= temp_mult_133(381);
partial_product_3(382) <= temp_mult_133(382);
partial_product_3(383) <= temp_mult_133(383);
partial_product_3(384) <= temp_mult_133(384);
partial_product_3(385) <= temp_mult_133(385);
partial_product_3(386) <= temp_mult_133(386);
partial_product_3(387) <= temp_mult_133(387);
partial_product_3(388) <= temp_mult_133(388);
partial_product_3(389) <= temp_mult_133(389);
partial_product_3(390) <= temp_mult_133(390);
partial_product_3(391) <= temp_mult_133(391);
partial_product_3(392) <= temp_mult_133(392);
partial_product_3(393) <= temp_mult_133(393);
partial_product_3(394) <= temp_mult_133(394);
partial_product_3(395) <= temp_mult_133(395);
partial_product_3(396) <= temp_mult_133(396);
partial_product_3(397) <= temp_mult_133(397);
partial_product_3(398) <= temp_mult_133(398);
partial_product_3(399) <= temp_mult_133(399);
partial_product_3(400) <= temp_mult_133(400);
partial_product_3(401) <= temp_mult_133(401);
partial_product_3(402) <= temp_mult_133(402);
partial_product_3(403) <= temp_mult_139(403);
partial_product_3(404) <= temp_mult_139(404);
partial_product_3(405) <= temp_mult_139(405);
partial_product_3(406) <= temp_mult_139(406);
partial_product_3(407) <= temp_mult_139(407);
partial_product_3(408) <= temp_mult_139(408);
partial_product_3(409) <= temp_mult_139(409);
partial_product_3(410) <= temp_mult_139(410);
partial_product_3(411) <= temp_mult_139(411);
partial_product_3(412) <= temp_mult_139(412);
partial_product_3(413) <= temp_mult_139(413);
partial_product_3(414) <= temp_mult_139(414);
partial_product_3(415) <= temp_mult_139(415);
partial_product_3(416) <= temp_mult_139(416);
partial_product_3(417) <= temp_mult_139(417);
partial_product_3(418) <= temp_mult_139(418);
partial_product_3(419) <= temp_mult_139(419);
partial_product_3(420) <= temp_mult_139(420);
partial_product_3(421) <= temp_mult_139(421);
partial_product_3(422) <= temp_mult_139(422);
partial_product_3(423) <= temp_mult_139(423);
partial_product_3(424) <= temp_mult_139(424);
partial_product_3(425) <= temp_mult_139(425);
partial_product_3(426) <= temp_mult_139(426);
partial_product_3(427) <= temp_mult_139(427);
partial_product_3(428) <= temp_mult_139(428);
partial_product_3(429) <= temp_mult_139(429);
partial_product_3(430) <= temp_mult_139(430);
partial_product_3(431) <= temp_mult_139(431);
partial_product_3(432) <= temp_mult_139(432);
partial_product_3(433) <= temp_mult_139(433);
partial_product_3(434) <= temp_mult_139(434);
partial_product_3(435) <= temp_mult_139(435);
partial_product_3(436) <= temp_mult_139(436);
partial_product_3(437) <= temp_mult_139(437);
partial_product_3(438) <= temp_mult_139(438);
partial_product_3(439) <= temp_mult_139(439);
partial_product_3(440) <= temp_mult_139(440);
partial_product_3(441) <= temp_mult_139(441);
partial_product_3(442) <= temp_mult_139(442);
partial_product_3(443) <= temp_mult_139(443);
partial_product_3(444) <= '0';
partial_product_3(445) <= '0';
partial_product_3(446) <= '0';
partial_product_3(447) <= temp_mult_158(447);
partial_product_3(448) <= temp_mult_158(448);
partial_product_3(449) <= temp_mult_158(449);
partial_product_3(450) <= temp_mult_158(450);
partial_product_3(451) <= temp_mult_158(451);
partial_product_3(452) <= temp_mult_158(452);
partial_product_3(453) <= temp_mult_158(453);
partial_product_3(454) <= temp_mult_158(454);
partial_product_3(455) <= temp_mult_158(455);
partial_product_3(456) <= temp_mult_158(456);
partial_product_3(457) <= temp_mult_158(457);
partial_product_3(458) <= temp_mult_158(458);
partial_product_3(459) <= temp_mult_158(459);
partial_product_3(460) <= temp_mult_158(460);
partial_product_3(461) <= temp_mult_158(461);
partial_product_3(462) <= temp_mult_158(462);
partial_product_3(463) <= temp_mult_158(463);
partial_product_3(464) <= temp_mult_158(464);
partial_product_3(465) <= temp_mult_158(465);
partial_product_3(466) <= temp_mult_158(466);
partial_product_3(467) <= temp_mult_158(467);
partial_product_3(468) <= temp_mult_158(468);
partial_product_3(469) <= temp_mult_158(469);
partial_product_3(470) <= temp_mult_158(470);
partial_product_3(471) <= temp_mult_158(471);
partial_product_3(472) <= temp_mult_158(472);
partial_product_3(473) <= temp_mult_158(473);
partial_product_3(474) <= temp_mult_158(474);
partial_product_3(475) <= temp_mult_158(475);
partial_product_3(476) <= temp_mult_158(476);
partial_product_3(477) <= temp_mult_158(477);
partial_product_3(478) <= temp_mult_158(478);
partial_product_3(479) <= temp_mult_158(479);
partial_product_3(480) <= temp_mult_158(480);
partial_product_3(481) <= temp_mult_158(481);
partial_product_3(482) <= temp_mult_158(482);
partial_product_3(483) <= temp_mult_158(483);
partial_product_3(484) <= temp_mult_158(484);
partial_product_3(485) <= temp_mult_158(485);
partial_product_3(486) <= temp_mult_158(486);
partial_product_3(487) <= temp_mult_158(487);
partial_product_3(488) <= '0';
partial_product_3(489) <= '0';
partial_product_3(490) <= '0';
partial_product_3(491) <= '0';
partial_product_3(492) <= '0';
partial_product_3(493) <= '0';
partial_product_3(494) <= '0';
partial_product_3(495) <= '0';
partial_product_3(496) <= '0';
partial_product_3(497) <= '0';
partial_product_3(498) <= '0';
partial_product_3(499) <= '0';
partial_product_3(500) <= '0';
partial_product_3(501) <= '0';
partial_product_3(502) <= '0';
partial_product_3(503) <= '0';
partial_product_3(504) <= '0';
partial_product_3(505) <= '0';
partial_product_3(506) <= '0';
partial_product_3(507) <= '0';
partial_product_3(508) <= '0';
partial_product_3(509) <= '0';
partial_product_3(510) <= '0';
partial_product_3(511) <= '0';
partial_product_3(512) <= '0';
partial_product_4(0) <= '0';
partial_product_4(1) <= '0';
partial_product_4(2) <= '0';
partial_product_4(3) <= '0';
partial_product_4(4) <= '0';
partial_product_4(5) <= '0';
partial_product_4(6) <= '0';
partial_product_4(7) <= '0';
partial_product_4(8) <= '0';
partial_product_4(9) <= '0';
partial_product_4(10) <= '0';
partial_product_4(11) <= '0';
partial_product_4(12) <= '0';
partial_product_4(13) <= '0';
partial_product_4(14) <= '0';
partial_product_4(15) <= '0';
partial_product_4(16) <= '0';
partial_product_4(17) <= '0';
partial_product_4(18) <= '0';
partial_product_4(19) <= '0';
partial_product_4(20) <= '0';
partial_product_4(21) <= '0';
partial_product_4(22) <= '0';
partial_product_4(23) <= '0';
partial_product_4(24) <= '0';
partial_product_4(25) <= '0';
partial_product_4(26) <= '0';
partial_product_4(27) <= '0';
partial_product_4(28) <= '0';
partial_product_4(29) <= '0';
partial_product_4(30) <= '0';
partial_product_4(31) <= '0';
partial_product_4(32) <= '0';
partial_product_4(33) <= '0';
partial_product_4(34) <= '0';
partial_product_4(35) <= '0';
partial_product_4(36) <= '0';
partial_product_4(37) <= '0';
partial_product_4(38) <= '0';
partial_product_4(39) <= '0';
partial_product_4(40) <= '0';
partial_product_4(41) <= '0';
partial_product_4(42) <= '0';
partial_product_4(43) <= '0';
partial_product_4(44) <= '0';
partial_product_4(45) <= '0';
partial_product_4(46) <= '0';
partial_product_4(47) <= '0';
partial_product_4(48) <= temp_mult_2(48);
partial_product_4(49) <= temp_mult_2(49);
partial_product_4(50) <= temp_mult_2(50);
partial_product_4(51) <= temp_mult_2(51);
partial_product_4(52) <= temp_mult_2(52);
partial_product_4(53) <= temp_mult_2(53);
partial_product_4(54) <= temp_mult_2(54);
partial_product_4(55) <= temp_mult_2(55);
partial_product_4(56) <= temp_mult_2(56);
partial_product_4(57) <= temp_mult_2(57);
partial_product_4(58) <= temp_mult_2(58);
partial_product_4(59) <= temp_mult_2(59);
partial_product_4(60) <= temp_mult_2(60);
partial_product_4(61) <= temp_mult_2(61);
partial_product_4(62) <= temp_mult_2(62);
partial_product_4(63) <= temp_mult_2(63);
partial_product_4(64) <= temp_mult_2(64);
partial_product_4(65) <= temp_mult_2(65);
partial_product_4(66) <= temp_mult_2(66);
partial_product_4(67) <= temp_mult_2(67);
partial_product_4(68) <= temp_mult_2(68);
partial_product_4(69) <= temp_mult_2(69);
partial_product_4(70) <= temp_mult_2(70);
partial_product_4(71) <= temp_mult_2(71);
partial_product_4(72) <= temp_mult_2(72);
partial_product_4(73) <= temp_mult_2(73);
partial_product_4(74) <= temp_mult_2(74);
partial_product_4(75) <= temp_mult_2(75);
partial_product_4(76) <= temp_mult_2(76);
partial_product_4(77) <= temp_mult_2(77);
partial_product_4(78) <= temp_mult_2(78);
partial_product_4(79) <= temp_mult_2(79);
partial_product_4(80) <= temp_mult_2(80);
partial_product_4(81) <= temp_mult_2(81);
partial_product_4(82) <= temp_mult_2(82);
partial_product_4(83) <= temp_mult_2(83);
partial_product_4(84) <= temp_mult_2(84);
partial_product_4(85) <= temp_mult_2(85);
partial_product_4(86) <= temp_mult_2(86);
partial_product_4(87) <= temp_mult_2(87);
partial_product_4(88) <= temp_mult_2(88);
partial_product_4(89) <= temp_mult_8(89);
partial_product_4(90) <= temp_mult_8(90);
partial_product_4(91) <= temp_mult_8(91);
partial_product_4(92) <= temp_mult_8(92);
partial_product_4(93) <= temp_mult_8(93);
partial_product_4(94) <= temp_mult_8(94);
partial_product_4(95) <= temp_mult_8(95);
partial_product_4(96) <= temp_mult_8(96);
partial_product_4(97) <= temp_mult_8(97);
partial_product_4(98) <= temp_mult_8(98);
partial_product_4(99) <= temp_mult_8(99);
partial_product_4(100) <= temp_mult_8(100);
partial_product_4(101) <= temp_mult_8(101);
partial_product_4(102) <= temp_mult_8(102);
partial_product_4(103) <= temp_mult_8(103);
partial_product_4(104) <= temp_mult_8(104);
partial_product_4(105) <= temp_mult_8(105);
partial_product_4(106) <= temp_mult_8(106);
partial_product_4(107) <= temp_mult_8(107);
partial_product_4(108) <= temp_mult_8(108);
partial_product_4(109) <= temp_mult_8(109);
partial_product_4(110) <= temp_mult_8(110);
partial_product_4(111) <= temp_mult_8(111);
partial_product_4(112) <= temp_mult_8(112);
partial_product_4(113) <= temp_mult_8(113);
partial_product_4(114) <= temp_mult_8(114);
partial_product_4(115) <= temp_mult_8(115);
partial_product_4(116) <= temp_mult_8(116);
partial_product_4(117) <= temp_mult_8(117);
partial_product_4(118) <= temp_mult_8(118);
partial_product_4(119) <= temp_mult_8(119);
partial_product_4(120) <= temp_mult_8(120);
partial_product_4(121) <= temp_mult_8(121);
partial_product_4(122) <= temp_mult_8(122);
partial_product_4(123) <= temp_mult_8(123);
partial_product_4(124) <= temp_mult_8(124);
partial_product_4(125) <= temp_mult_8(125);
partial_product_4(126) <= temp_mult_8(126);
partial_product_4(127) <= temp_mult_8(127);
partial_product_4(128) <= temp_mult_8(128);
partial_product_4(129) <= temp_mult_8(129);
partial_product_4(130) <= temp_mult_14(130);
partial_product_4(131) <= temp_mult_14(131);
partial_product_4(132) <= temp_mult_14(132);
partial_product_4(133) <= temp_mult_14(133);
partial_product_4(134) <= temp_mult_14(134);
partial_product_4(135) <= temp_mult_14(135);
partial_product_4(136) <= temp_mult_14(136);
partial_product_4(137) <= temp_mult_14(137);
partial_product_4(138) <= temp_mult_14(138);
partial_product_4(139) <= temp_mult_14(139);
partial_product_4(140) <= temp_mult_14(140);
partial_product_4(141) <= temp_mult_14(141);
partial_product_4(142) <= temp_mult_14(142);
partial_product_4(143) <= temp_mult_14(143);
partial_product_4(144) <= temp_mult_14(144);
partial_product_4(145) <= temp_mult_14(145);
partial_product_4(146) <= temp_mult_14(146);
partial_product_4(147) <= temp_mult_14(147);
partial_product_4(148) <= temp_mult_14(148);
partial_product_4(149) <= temp_mult_14(149);
partial_product_4(150) <= temp_mult_14(150);
partial_product_4(151) <= temp_mult_14(151);
partial_product_4(152) <= temp_mult_14(152);
partial_product_4(153) <= temp_mult_14(153);
partial_product_4(154) <= temp_mult_14(154);
partial_product_4(155) <= temp_mult_14(155);
partial_product_4(156) <= temp_mult_14(156);
partial_product_4(157) <= temp_mult_14(157);
partial_product_4(158) <= temp_mult_14(158);
partial_product_4(159) <= temp_mult_14(159);
partial_product_4(160) <= temp_mult_14(160);
partial_product_4(161) <= temp_mult_14(161);
partial_product_4(162) <= temp_mult_14(162);
partial_product_4(163) <= temp_mult_14(163);
partial_product_4(164) <= temp_mult_14(164);
partial_product_4(165) <= temp_mult_14(165);
partial_product_4(166) <= temp_mult_14(166);
partial_product_4(167) <= temp_mult_14(167);
partial_product_4(168) <= temp_mult_14(168);
partial_product_4(169) <= temp_mult_14(169);
partial_product_4(170) <= temp_mult_14(170);
partial_product_4(171) <= temp_mult_43(171);
partial_product_4(172) <= temp_mult_43(172);
partial_product_4(173) <= temp_mult_43(173);
partial_product_4(174) <= temp_mult_43(174);
partial_product_4(175) <= temp_mult_43(175);
partial_product_4(176) <= temp_mult_43(176);
partial_product_4(177) <= temp_mult_43(177);
partial_product_4(178) <= temp_mult_43(178);
partial_product_4(179) <= temp_mult_43(179);
partial_product_4(180) <= temp_mult_43(180);
partial_product_4(181) <= temp_mult_43(181);
partial_product_4(182) <= temp_mult_43(182);
partial_product_4(183) <= temp_mult_43(183);
partial_product_4(184) <= temp_mult_43(184);
partial_product_4(185) <= temp_mult_43(185);
partial_product_4(186) <= temp_mult_43(186);
partial_product_4(187) <= temp_mult_43(187);
partial_product_4(188) <= temp_mult_43(188);
partial_product_4(189) <= temp_mult_43(189);
partial_product_4(190) <= temp_mult_43(190);
partial_product_4(191) <= temp_mult_43(191);
partial_product_4(192) <= temp_mult_43(192);
partial_product_4(193) <= temp_mult_43(193);
partial_product_4(194) <= temp_mult_43(194);
partial_product_4(195) <= temp_mult_43(195);
partial_product_4(196) <= temp_mult_43(196);
partial_product_4(197) <= temp_mult_43(197);
partial_product_4(198) <= temp_mult_43(198);
partial_product_4(199) <= temp_mult_43(199);
partial_product_4(200) <= temp_mult_43(200);
partial_product_4(201) <= temp_mult_43(201);
partial_product_4(202) <= temp_mult_43(202);
partial_product_4(203) <= temp_mult_43(203);
partial_product_4(204) <= temp_mult_43(204);
partial_product_4(205) <= temp_mult_43(205);
partial_product_4(206) <= temp_mult_43(206);
partial_product_4(207) <= temp_mult_43(207);
partial_product_4(208) <= temp_mult_43(208);
partial_product_4(209) <= temp_mult_43(209);
partial_product_4(210) <= temp_mult_43(210);
partial_product_4(211) <= temp_mult_43(211);
partial_product_4(212) <= temp_mult_52(212);
partial_product_4(213) <= temp_mult_52(213);
partial_product_4(214) <= temp_mult_52(214);
partial_product_4(215) <= temp_mult_52(215);
partial_product_4(216) <= temp_mult_52(216);
partial_product_4(217) <= temp_mult_52(217);
partial_product_4(218) <= temp_mult_52(218);
partial_product_4(219) <= temp_mult_52(219);
partial_product_4(220) <= temp_mult_52(220);
partial_product_4(221) <= temp_mult_52(221);
partial_product_4(222) <= temp_mult_52(222);
partial_product_4(223) <= temp_mult_52(223);
partial_product_4(224) <= temp_mult_52(224);
partial_product_4(225) <= temp_mult_52(225);
partial_product_4(226) <= temp_mult_52(226);
partial_product_4(227) <= temp_mult_52(227);
partial_product_4(228) <= temp_mult_52(228);
partial_product_4(229) <= temp_mult_52(229);
partial_product_4(230) <= temp_mult_52(230);
partial_product_4(231) <= temp_mult_52(231);
partial_product_4(232) <= temp_mult_52(232);
partial_product_4(233) <= temp_mult_52(233);
partial_product_4(234) <= temp_mult_52(234);
partial_product_4(235) <= temp_mult_52(235);
partial_product_4(236) <= temp_mult_52(236);
partial_product_4(237) <= temp_mult_52(237);
partial_product_4(238) <= temp_mult_52(238);
partial_product_4(239) <= temp_mult_52(239);
partial_product_4(240) <= temp_mult_52(240);
partial_product_4(241) <= temp_mult_52(241);
partial_product_4(242) <= temp_mult_52(242);
partial_product_4(243) <= temp_mult_52(243);
partial_product_4(244) <= temp_mult_52(244);
partial_product_4(245) <= temp_mult_52(245);
partial_product_4(246) <= temp_mult_52(246);
partial_product_4(247) <= temp_mult_52(247);
partial_product_4(248) <= temp_mult_52(248);
partial_product_4(249) <= temp_mult_52(249);
partial_product_4(250) <= temp_mult_52(250);
partial_product_4(251) <= temp_mult_52(251);
partial_product_4(252) <= temp_mult_52(252);
partial_product_4(253) <= temp_mult_61(253);
partial_product_4(254) <= temp_mult_61(254);
partial_product_4(255) <= temp_mult_61(255);
partial_product_4(256) <= temp_mult_61(256);
partial_product_4(257) <= temp_mult_61(257);
partial_product_4(258) <= temp_mult_61(258);
partial_product_4(259) <= temp_mult_61(259);
partial_product_4(260) <= temp_mult_61(260);
partial_product_4(261) <= temp_mult_61(261);
partial_product_4(262) <= temp_mult_61(262);
partial_product_4(263) <= temp_mult_61(263);
partial_product_4(264) <= temp_mult_61(264);
partial_product_4(265) <= temp_mult_61(265);
partial_product_4(266) <= temp_mult_61(266);
partial_product_4(267) <= temp_mult_61(267);
partial_product_4(268) <= temp_mult_61(268);
partial_product_4(269) <= temp_mult_61(269);
partial_product_4(270) <= temp_mult_61(270);
partial_product_4(271) <= temp_mult_61(271);
partial_product_4(272) <= temp_mult_61(272);
partial_product_4(273) <= temp_mult_61(273);
partial_product_4(274) <= temp_mult_61(274);
partial_product_4(275) <= temp_mult_61(275);
partial_product_4(276) <= temp_mult_61(276);
partial_product_4(277) <= temp_mult_61(277);
partial_product_4(278) <= temp_mult_61(278);
partial_product_4(279) <= temp_mult_61(279);
partial_product_4(280) <= temp_mult_61(280);
partial_product_4(281) <= temp_mult_61(281);
partial_product_4(282) <= temp_mult_61(282);
partial_product_4(283) <= temp_mult_61(283);
partial_product_4(284) <= temp_mult_61(284);
partial_product_4(285) <= temp_mult_61(285);
partial_product_4(286) <= temp_mult_61(286);
partial_product_4(287) <= temp_mult_61(287);
partial_product_4(288) <= temp_mult_61(288);
partial_product_4(289) <= temp_mult_61(289);
partial_product_4(290) <= temp_mult_61(290);
partial_product_4(291) <= temp_mult_61(291);
partial_product_4(292) <= temp_mult_61(292);
partial_product_4(293) <= temp_mult_61(293);
partial_product_4(294) <= temp_mult_70(294);
partial_product_4(295) <= temp_mult_70(295);
partial_product_4(296) <= temp_mult_70(296);
partial_product_4(297) <= temp_mult_70(297);
partial_product_4(298) <= temp_mult_70(298);
partial_product_4(299) <= temp_mult_70(299);
partial_product_4(300) <= temp_mult_70(300);
partial_product_4(301) <= temp_mult_70(301);
partial_product_4(302) <= temp_mult_70(302);
partial_product_4(303) <= temp_mult_70(303);
partial_product_4(304) <= temp_mult_70(304);
partial_product_4(305) <= temp_mult_70(305);
partial_product_4(306) <= temp_mult_70(306);
partial_product_4(307) <= temp_mult_70(307);
partial_product_4(308) <= temp_mult_70(308);
partial_product_4(309) <= temp_mult_70(309);
partial_product_4(310) <= temp_mult_70(310);
partial_product_4(311) <= temp_mult_70(311);
partial_product_4(312) <= temp_mult_70(312);
partial_product_4(313) <= temp_mult_70(313);
partial_product_4(314) <= temp_mult_70(314);
partial_product_4(315) <= temp_mult_70(315);
partial_product_4(316) <= temp_mult_70(316);
partial_product_4(317) <= temp_mult_70(317);
partial_product_4(318) <= temp_mult_70(318);
partial_product_4(319) <= temp_mult_70(319);
partial_product_4(320) <= temp_mult_70(320);
partial_product_4(321) <= temp_mult_70(321);
partial_product_4(322) <= temp_mult_70(322);
partial_product_4(323) <= temp_mult_70(323);
partial_product_4(324) <= temp_mult_70(324);
partial_product_4(325) <= temp_mult_70(325);
partial_product_4(326) <= temp_mult_70(326);
partial_product_4(327) <= temp_mult_70(327);
partial_product_4(328) <= temp_mult_70(328);
partial_product_4(329) <= temp_mult_70(329);
partial_product_4(330) <= temp_mult_70(330);
partial_product_4(331) <= temp_mult_70(331);
partial_product_4(332) <= temp_mult_70(332);
partial_product_4(333) <= temp_mult_70(333);
partial_product_4(334) <= temp_mult_70(334);
partial_product_4(335) <= temp_mult_79(335);
partial_product_4(336) <= temp_mult_79(336);
partial_product_4(337) <= temp_mult_79(337);
partial_product_4(338) <= temp_mult_79(338);
partial_product_4(339) <= temp_mult_79(339);
partial_product_4(340) <= temp_mult_79(340);
partial_product_4(341) <= temp_mult_79(341);
partial_product_4(342) <= temp_mult_79(342);
partial_product_4(343) <= temp_mult_79(343);
partial_product_4(344) <= temp_mult_79(344);
partial_product_4(345) <= temp_mult_79(345);
partial_product_4(346) <= temp_mult_79(346);
partial_product_4(347) <= temp_mult_79(347);
partial_product_4(348) <= temp_mult_79(348);
partial_product_4(349) <= temp_mult_79(349);
partial_product_4(350) <= temp_mult_79(350);
partial_product_4(351) <= temp_mult_79(351);
partial_product_4(352) <= temp_mult_79(352);
partial_product_4(353) <= temp_mult_79(353);
partial_product_4(354) <= temp_mult_79(354);
partial_product_4(355) <= temp_mult_79(355);
partial_product_4(356) <= temp_mult_79(356);
partial_product_4(357) <= temp_mult_79(357);
partial_product_4(358) <= temp_mult_79(358);
partial_product_4(359) <= temp_mult_79(359);
partial_product_4(360) <= temp_mult_79(360);
partial_product_4(361) <= temp_mult_79(361);
partial_product_4(362) <= temp_mult_79(362);
partial_product_4(363) <= temp_mult_79(363);
partial_product_4(364) <= temp_mult_79(364);
partial_product_4(365) <= temp_mult_79(365);
partial_product_4(366) <= temp_mult_79(366);
partial_product_4(367) <= temp_mult_79(367);
partial_product_4(368) <= temp_mult_79(368);
partial_product_4(369) <= temp_mult_79(369);
partial_product_4(370) <= temp_mult_79(370);
partial_product_4(371) <= temp_mult_79(371);
partial_product_4(372) <= temp_mult_79(372);
partial_product_4(373) <= temp_mult_79(373);
partial_product_4(374) <= temp_mult_79(374);
partial_product_4(375) <= temp_mult_79(375);
partial_product_4(376) <= '0';
partial_product_4(377) <= '0';
partial_product_4(378) <= '0';
partial_product_4(379) <= temp_mult_138(379);
partial_product_4(380) <= temp_mult_138(380);
partial_product_4(381) <= temp_mult_138(381);
partial_product_4(382) <= temp_mult_138(382);
partial_product_4(383) <= temp_mult_138(383);
partial_product_4(384) <= temp_mult_138(384);
partial_product_4(385) <= temp_mult_138(385);
partial_product_4(386) <= temp_mult_138(386);
partial_product_4(387) <= temp_mult_138(387);
partial_product_4(388) <= temp_mult_138(388);
partial_product_4(389) <= temp_mult_138(389);
partial_product_4(390) <= temp_mult_138(390);
partial_product_4(391) <= temp_mult_138(391);
partial_product_4(392) <= temp_mult_138(392);
partial_product_4(393) <= temp_mult_138(393);
partial_product_4(394) <= temp_mult_138(394);
partial_product_4(395) <= temp_mult_138(395);
partial_product_4(396) <= temp_mult_138(396);
partial_product_4(397) <= temp_mult_138(397);
partial_product_4(398) <= temp_mult_138(398);
partial_product_4(399) <= temp_mult_138(399);
partial_product_4(400) <= temp_mult_138(400);
partial_product_4(401) <= temp_mult_138(401);
partial_product_4(402) <= temp_mult_138(402);
partial_product_4(403) <= temp_mult_138(403);
partial_product_4(404) <= temp_mult_138(404);
partial_product_4(405) <= temp_mult_138(405);
partial_product_4(406) <= temp_mult_138(406);
partial_product_4(407) <= temp_mult_138(407);
partial_product_4(408) <= temp_mult_138(408);
partial_product_4(409) <= temp_mult_138(409);
partial_product_4(410) <= temp_mult_138(410);
partial_product_4(411) <= temp_mult_138(411);
partial_product_4(412) <= temp_mult_138(412);
partial_product_4(413) <= temp_mult_138(413);
partial_product_4(414) <= temp_mult_138(414);
partial_product_4(415) <= temp_mult_138(415);
partial_product_4(416) <= temp_mult_138(416);
partial_product_4(417) <= temp_mult_138(417);
partial_product_4(418) <= temp_mult_138(418);
partial_product_4(419) <= temp_mult_138(419);
partial_product_4(420) <= temp_mult_144(420);
partial_product_4(421) <= temp_mult_144(421);
partial_product_4(422) <= temp_mult_144(422);
partial_product_4(423) <= temp_mult_144(423);
partial_product_4(424) <= temp_mult_144(424);
partial_product_4(425) <= temp_mult_144(425);
partial_product_4(426) <= temp_mult_144(426);
partial_product_4(427) <= temp_mult_144(427);
partial_product_4(428) <= temp_mult_144(428);
partial_product_4(429) <= temp_mult_144(429);
partial_product_4(430) <= temp_mult_144(430);
partial_product_4(431) <= temp_mult_144(431);
partial_product_4(432) <= temp_mult_144(432);
partial_product_4(433) <= temp_mult_144(433);
partial_product_4(434) <= temp_mult_144(434);
partial_product_4(435) <= temp_mult_144(435);
partial_product_4(436) <= temp_mult_144(436);
partial_product_4(437) <= temp_mult_144(437);
partial_product_4(438) <= temp_mult_144(438);
partial_product_4(439) <= temp_mult_144(439);
partial_product_4(440) <= temp_mult_144(440);
partial_product_4(441) <= temp_mult_144(441);
partial_product_4(442) <= temp_mult_144(442);
partial_product_4(443) <= temp_mult_144(443);
partial_product_4(444) <= temp_mult_144(444);
partial_product_4(445) <= temp_mult_144(445);
partial_product_4(446) <= temp_mult_144(446);
partial_product_4(447) <= temp_mult_144(447);
partial_product_4(448) <= temp_mult_144(448);
partial_product_4(449) <= temp_mult_144(449);
partial_product_4(450) <= temp_mult_144(450);
partial_product_4(451) <= temp_mult_144(451);
partial_product_4(452) <= temp_mult_144(452);
partial_product_4(453) <= temp_mult_144(453);
partial_product_4(454) <= temp_mult_144(454);
partial_product_4(455) <= temp_mult_144(455);
partial_product_4(456) <= temp_mult_144(456);
partial_product_4(457) <= temp_mult_144(457);
partial_product_4(458) <= temp_mult_144(458);
partial_product_4(459) <= temp_mult_144(459);
partial_product_4(460) <= temp_mult_144(460);
partial_product_4(461) <= '0';
partial_product_4(462) <= '0';
partial_product_4(463) <= '0';
partial_product_4(464) <= '0';
partial_product_4(465) <= '0';
partial_product_4(466) <= '0';
partial_product_4(467) <= '0';
partial_product_4(468) <= '0';
partial_product_4(469) <= '0';
partial_product_4(470) <= '0';
partial_product_4(471) <= '0';
partial_product_4(472) <= '0';
partial_product_4(473) <= '0';
partial_product_4(474) <= '0';
partial_product_4(475) <= '0';
partial_product_4(476) <= '0';
partial_product_4(477) <= '0';
partial_product_4(478) <= '0';
partial_product_4(479) <= '0';
partial_product_4(480) <= '0';
partial_product_4(481) <= '0';
partial_product_4(482) <= '0';
partial_product_4(483) <= '0';
partial_product_4(484) <= '0';
partial_product_4(485) <= '0';
partial_product_4(486) <= '0';
partial_product_4(487) <= '0';
partial_product_4(488) <= '0';
partial_product_4(489) <= '0';
partial_product_4(490) <= '0';
partial_product_4(491) <= '0';
partial_product_4(492) <= '0';
partial_product_4(493) <= '0';
partial_product_4(494) <= '0';
partial_product_4(495) <= '0';
partial_product_4(496) <= '0';
partial_product_4(497) <= '0';
partial_product_4(498) <= '0';
partial_product_4(499) <= '0';
partial_product_4(500) <= '0';
partial_product_4(501) <= '0';
partial_product_4(502) <= '0';
partial_product_4(503) <= '0';
partial_product_4(504) <= '0';
partial_product_4(505) <= '0';
partial_product_4(506) <= '0';
partial_product_4(507) <= '0';
partial_product_4(508) <= '0';
partial_product_4(509) <= '0';
partial_product_4(510) <= '0';
partial_product_4(511) <= '0';
partial_product_4(512) <= '0';
partial_product_5(0) <= '0';
partial_product_5(1) <= '0';
partial_product_5(2) <= '0';
partial_product_5(3) <= '0';
partial_product_5(4) <= '0';
partial_product_5(5) <= '0';
partial_product_5(6) <= '0';
partial_product_5(7) <= '0';
partial_product_5(8) <= '0';
partial_product_5(9) <= '0';
partial_product_5(10) <= '0';
partial_product_5(11) <= '0';
partial_product_5(12) <= '0';
partial_product_5(13) <= '0';
partial_product_5(14) <= '0';
partial_product_5(15) <= '0';
partial_product_5(16) <= '0';
partial_product_5(17) <= '0';
partial_product_5(18) <= '0';
partial_product_5(19) <= '0';
partial_product_5(20) <= '0';
partial_product_5(21) <= '0';
partial_product_5(22) <= '0';
partial_product_5(23) <= '0';
partial_product_5(24) <= '0';
partial_product_5(25) <= '0';
partial_product_5(26) <= '0';
partial_product_5(27) <= '0';
partial_product_5(28) <= '0';
partial_product_5(29) <= '0';
partial_product_5(30) <= '0';
partial_product_5(31) <= '0';
partial_product_5(32) <= '0';
partial_product_5(33) <= '0';
partial_product_5(34) <= '0';
partial_product_5(35) <= '0';
partial_product_5(36) <= '0';
partial_product_5(37) <= '0';
partial_product_5(38) <= '0';
partial_product_5(39) <= '0';
partial_product_5(40) <= '0';
partial_product_5(41) <= '0';
partial_product_5(42) <= '0';
partial_product_5(43) <= '0';
partial_product_5(44) <= '0';
partial_product_5(45) <= '0';
partial_product_5(46) <= '0';
partial_product_5(47) <= '0';
partial_product_5(48) <= '0';
partial_product_5(49) <= '0';
partial_product_5(50) <= '0';
partial_product_5(51) <= temp_mult_15(51);
partial_product_5(52) <= temp_mult_15(52);
partial_product_5(53) <= temp_mult_15(53);
partial_product_5(54) <= temp_mult_15(54);
partial_product_5(55) <= temp_mult_15(55);
partial_product_5(56) <= temp_mult_15(56);
partial_product_5(57) <= temp_mult_15(57);
partial_product_5(58) <= temp_mult_15(58);
partial_product_5(59) <= temp_mult_15(59);
partial_product_5(60) <= temp_mult_15(60);
partial_product_5(61) <= temp_mult_15(61);
partial_product_5(62) <= temp_mult_15(62);
partial_product_5(63) <= temp_mult_15(63);
partial_product_5(64) <= temp_mult_15(64);
partial_product_5(65) <= temp_mult_15(65);
partial_product_5(66) <= temp_mult_15(66);
partial_product_5(67) <= temp_mult_15(67);
partial_product_5(68) <= temp_mult_15(68);
partial_product_5(69) <= temp_mult_15(69);
partial_product_5(70) <= temp_mult_15(70);
partial_product_5(71) <= temp_mult_15(71);
partial_product_5(72) <= temp_mult_15(72);
partial_product_5(73) <= temp_mult_15(73);
partial_product_5(74) <= temp_mult_15(74);
partial_product_5(75) <= temp_mult_15(75);
partial_product_5(76) <= temp_mult_15(76);
partial_product_5(77) <= temp_mult_15(77);
partial_product_5(78) <= temp_mult_15(78);
partial_product_5(79) <= temp_mult_15(79);
partial_product_5(80) <= temp_mult_15(80);
partial_product_5(81) <= temp_mult_15(81);
partial_product_5(82) <= temp_mult_15(82);
partial_product_5(83) <= temp_mult_15(83);
partial_product_5(84) <= temp_mult_15(84);
partial_product_5(85) <= temp_mult_15(85);
partial_product_5(86) <= temp_mult_15(86);
partial_product_5(87) <= temp_mult_15(87);
partial_product_5(88) <= temp_mult_15(88);
partial_product_5(89) <= temp_mult_15(89);
partial_product_5(90) <= temp_mult_15(90);
partial_product_5(91) <= temp_mult_15(91);
partial_product_5(92) <= temp_mult_21(92);
partial_product_5(93) <= temp_mult_21(93);
partial_product_5(94) <= temp_mult_21(94);
partial_product_5(95) <= temp_mult_21(95);
partial_product_5(96) <= temp_mult_21(96);
partial_product_5(97) <= temp_mult_21(97);
partial_product_5(98) <= temp_mult_21(98);
partial_product_5(99) <= temp_mult_21(99);
partial_product_5(100) <= temp_mult_21(100);
partial_product_5(101) <= temp_mult_21(101);
partial_product_5(102) <= temp_mult_21(102);
partial_product_5(103) <= temp_mult_21(103);
partial_product_5(104) <= temp_mult_21(104);
partial_product_5(105) <= temp_mult_21(105);
partial_product_5(106) <= temp_mult_21(106);
partial_product_5(107) <= temp_mult_21(107);
partial_product_5(108) <= temp_mult_21(108);
partial_product_5(109) <= temp_mult_21(109);
partial_product_5(110) <= temp_mult_21(110);
partial_product_5(111) <= temp_mult_21(111);
partial_product_5(112) <= temp_mult_21(112);
partial_product_5(113) <= temp_mult_21(113);
partial_product_5(114) <= temp_mult_21(114);
partial_product_5(115) <= temp_mult_21(115);
partial_product_5(116) <= temp_mult_21(116);
partial_product_5(117) <= temp_mult_21(117);
partial_product_5(118) <= temp_mult_21(118);
partial_product_5(119) <= temp_mult_21(119);
partial_product_5(120) <= temp_mult_21(120);
partial_product_5(121) <= temp_mult_21(121);
partial_product_5(122) <= temp_mult_21(122);
partial_product_5(123) <= temp_mult_21(123);
partial_product_5(124) <= temp_mult_21(124);
partial_product_5(125) <= temp_mult_21(125);
partial_product_5(126) <= temp_mult_21(126);
partial_product_5(127) <= temp_mult_21(127);
partial_product_5(128) <= temp_mult_21(128);
partial_product_5(129) <= temp_mult_21(129);
partial_product_5(130) <= temp_mult_21(130);
partial_product_5(131) <= temp_mult_21(131);
partial_product_5(132) <= temp_mult_21(132);
partial_product_5(133) <= temp_mult_27(133);
partial_product_5(134) <= temp_mult_27(134);
partial_product_5(135) <= temp_mult_27(135);
partial_product_5(136) <= temp_mult_27(136);
partial_product_5(137) <= temp_mult_27(137);
partial_product_5(138) <= temp_mult_27(138);
partial_product_5(139) <= temp_mult_27(139);
partial_product_5(140) <= temp_mult_27(140);
partial_product_5(141) <= temp_mult_27(141);
partial_product_5(142) <= temp_mult_27(142);
partial_product_5(143) <= temp_mult_27(143);
partial_product_5(144) <= temp_mult_27(144);
partial_product_5(145) <= temp_mult_27(145);
partial_product_5(146) <= temp_mult_27(146);
partial_product_5(147) <= temp_mult_27(147);
partial_product_5(148) <= temp_mult_27(148);
partial_product_5(149) <= temp_mult_27(149);
partial_product_5(150) <= temp_mult_27(150);
partial_product_5(151) <= temp_mult_27(151);
partial_product_5(152) <= temp_mult_27(152);
partial_product_5(153) <= temp_mult_27(153);
partial_product_5(154) <= temp_mult_27(154);
partial_product_5(155) <= temp_mult_27(155);
partial_product_5(156) <= temp_mult_27(156);
partial_product_5(157) <= temp_mult_27(157);
partial_product_5(158) <= temp_mult_27(158);
partial_product_5(159) <= temp_mult_27(159);
partial_product_5(160) <= temp_mult_27(160);
partial_product_5(161) <= temp_mult_27(161);
partial_product_5(162) <= temp_mult_27(162);
partial_product_5(163) <= temp_mult_27(163);
partial_product_5(164) <= temp_mult_27(164);
partial_product_5(165) <= temp_mult_27(165);
partial_product_5(166) <= temp_mult_27(166);
partial_product_5(167) <= temp_mult_27(167);
partial_product_5(168) <= temp_mult_27(168);
partial_product_5(169) <= temp_mult_27(169);
partial_product_5(170) <= temp_mult_27(170);
partial_product_5(171) <= temp_mult_27(171);
partial_product_5(172) <= temp_mult_27(172);
partial_product_5(173) <= temp_mult_27(173);
partial_product_5(174) <= temp_mult_33(174);
partial_product_5(175) <= temp_mult_33(175);
partial_product_5(176) <= temp_mult_33(176);
partial_product_5(177) <= temp_mult_33(177);
partial_product_5(178) <= temp_mult_33(178);
partial_product_5(179) <= temp_mult_33(179);
partial_product_5(180) <= temp_mult_33(180);
partial_product_5(181) <= temp_mult_33(181);
partial_product_5(182) <= temp_mult_33(182);
partial_product_5(183) <= temp_mult_33(183);
partial_product_5(184) <= temp_mult_33(184);
partial_product_5(185) <= temp_mult_33(185);
partial_product_5(186) <= temp_mult_33(186);
partial_product_5(187) <= temp_mult_33(187);
partial_product_5(188) <= temp_mult_33(188);
partial_product_5(189) <= temp_mult_33(189);
partial_product_5(190) <= temp_mult_33(190);
partial_product_5(191) <= temp_mult_33(191);
partial_product_5(192) <= temp_mult_33(192);
partial_product_5(193) <= temp_mult_33(193);
partial_product_5(194) <= temp_mult_33(194);
partial_product_5(195) <= temp_mult_33(195);
partial_product_5(196) <= temp_mult_33(196);
partial_product_5(197) <= temp_mult_33(197);
partial_product_5(198) <= temp_mult_33(198);
partial_product_5(199) <= temp_mult_33(199);
partial_product_5(200) <= temp_mult_33(200);
partial_product_5(201) <= temp_mult_33(201);
partial_product_5(202) <= temp_mult_33(202);
partial_product_5(203) <= temp_mult_33(203);
partial_product_5(204) <= temp_mult_33(204);
partial_product_5(205) <= temp_mult_33(205);
partial_product_5(206) <= temp_mult_33(206);
partial_product_5(207) <= temp_mult_33(207);
partial_product_5(208) <= temp_mult_33(208);
partial_product_5(209) <= temp_mult_33(209);
partial_product_5(210) <= temp_mult_33(210);
partial_product_5(211) <= temp_mult_33(211);
partial_product_5(212) <= temp_mult_33(212);
partial_product_5(213) <= temp_mult_33(213);
partial_product_5(214) <= temp_mult_33(214);
partial_product_5(215) <= temp_mult_39(215);
partial_product_5(216) <= temp_mult_39(216);
partial_product_5(217) <= temp_mult_39(217);
partial_product_5(218) <= temp_mult_39(218);
partial_product_5(219) <= temp_mult_39(219);
partial_product_5(220) <= temp_mult_39(220);
partial_product_5(221) <= temp_mult_39(221);
partial_product_5(222) <= temp_mult_39(222);
partial_product_5(223) <= temp_mult_39(223);
partial_product_5(224) <= temp_mult_39(224);
partial_product_5(225) <= temp_mult_39(225);
partial_product_5(226) <= temp_mult_39(226);
partial_product_5(227) <= temp_mult_39(227);
partial_product_5(228) <= temp_mult_39(228);
partial_product_5(229) <= temp_mult_39(229);
partial_product_5(230) <= temp_mult_39(230);
partial_product_5(231) <= temp_mult_39(231);
partial_product_5(232) <= temp_mult_39(232);
partial_product_5(233) <= temp_mult_39(233);
partial_product_5(234) <= temp_mult_39(234);
partial_product_5(235) <= temp_mult_39(235);
partial_product_5(236) <= temp_mult_39(236);
partial_product_5(237) <= temp_mult_39(237);
partial_product_5(238) <= temp_mult_39(238);
partial_product_5(239) <= temp_mult_39(239);
partial_product_5(240) <= temp_mult_39(240);
partial_product_5(241) <= temp_mult_39(241);
partial_product_5(242) <= temp_mult_39(242);
partial_product_5(243) <= temp_mult_39(243);
partial_product_5(244) <= temp_mult_39(244);
partial_product_5(245) <= temp_mult_39(245);
partial_product_5(246) <= temp_mult_39(246);
partial_product_5(247) <= temp_mult_39(247);
partial_product_5(248) <= temp_mult_39(248);
partial_product_5(249) <= temp_mult_39(249);
partial_product_5(250) <= temp_mult_39(250);
partial_product_5(251) <= temp_mult_39(251);
partial_product_5(252) <= temp_mult_39(252);
partial_product_5(253) <= temp_mult_39(253);
partial_product_5(254) <= temp_mult_39(254);
partial_product_5(255) <= temp_mult_39(255);
partial_product_5(256) <= temp_mult_120(256);
partial_product_5(257) <= temp_mult_120(257);
partial_product_5(258) <= temp_mult_120(258);
partial_product_5(259) <= temp_mult_120(259);
partial_product_5(260) <= temp_mult_120(260);
partial_product_5(261) <= temp_mult_120(261);
partial_product_5(262) <= temp_mult_120(262);
partial_product_5(263) <= temp_mult_120(263);
partial_product_5(264) <= temp_mult_120(264);
partial_product_5(265) <= temp_mult_120(265);
partial_product_5(266) <= temp_mult_120(266);
partial_product_5(267) <= temp_mult_120(267);
partial_product_5(268) <= temp_mult_120(268);
partial_product_5(269) <= temp_mult_120(269);
partial_product_5(270) <= temp_mult_120(270);
partial_product_5(271) <= temp_mult_120(271);
partial_product_5(272) <= temp_mult_120(272);
partial_product_5(273) <= temp_mult_120(273);
partial_product_5(274) <= temp_mult_120(274);
partial_product_5(275) <= temp_mult_120(275);
partial_product_5(276) <= temp_mult_120(276);
partial_product_5(277) <= temp_mult_120(277);
partial_product_5(278) <= temp_mult_120(278);
partial_product_5(279) <= temp_mult_120(279);
partial_product_5(280) <= temp_mult_120(280);
partial_product_5(281) <= temp_mult_120(281);
partial_product_5(282) <= temp_mult_120(282);
partial_product_5(283) <= temp_mult_120(283);
partial_product_5(284) <= temp_mult_120(284);
partial_product_5(285) <= temp_mult_120(285);
partial_product_5(286) <= temp_mult_120(286);
partial_product_5(287) <= temp_mult_120(287);
partial_product_5(288) <= temp_mult_120(288);
partial_product_5(289) <= temp_mult_120(289);
partial_product_5(290) <= temp_mult_120(290);
partial_product_5(291) <= temp_mult_120(291);
partial_product_5(292) <= temp_mult_120(292);
partial_product_5(293) <= temp_mult_120(293);
partial_product_5(294) <= temp_mult_120(294);
partial_product_5(295) <= temp_mult_120(295);
partial_product_5(296) <= temp_mult_120(296);
partial_product_5(297) <= temp_mult_126(297);
partial_product_5(298) <= temp_mult_126(298);
partial_product_5(299) <= temp_mult_126(299);
partial_product_5(300) <= temp_mult_126(300);
partial_product_5(301) <= temp_mult_126(301);
partial_product_5(302) <= temp_mult_126(302);
partial_product_5(303) <= temp_mult_126(303);
partial_product_5(304) <= temp_mult_126(304);
partial_product_5(305) <= temp_mult_126(305);
partial_product_5(306) <= temp_mult_126(306);
partial_product_5(307) <= temp_mult_126(307);
partial_product_5(308) <= temp_mult_126(308);
partial_product_5(309) <= temp_mult_126(309);
partial_product_5(310) <= temp_mult_126(310);
partial_product_5(311) <= temp_mult_126(311);
partial_product_5(312) <= temp_mult_126(312);
partial_product_5(313) <= temp_mult_126(313);
partial_product_5(314) <= temp_mult_126(314);
partial_product_5(315) <= temp_mult_126(315);
partial_product_5(316) <= temp_mult_126(316);
partial_product_5(317) <= temp_mult_126(317);
partial_product_5(318) <= temp_mult_126(318);
partial_product_5(319) <= temp_mult_126(319);
partial_product_5(320) <= temp_mult_126(320);
partial_product_5(321) <= temp_mult_126(321);
partial_product_5(322) <= temp_mult_126(322);
partial_product_5(323) <= temp_mult_126(323);
partial_product_5(324) <= temp_mult_126(324);
partial_product_5(325) <= temp_mult_126(325);
partial_product_5(326) <= temp_mult_126(326);
partial_product_5(327) <= temp_mult_126(327);
partial_product_5(328) <= temp_mult_126(328);
partial_product_5(329) <= temp_mult_126(329);
partial_product_5(330) <= temp_mult_126(330);
partial_product_5(331) <= temp_mult_126(331);
partial_product_5(332) <= temp_mult_126(332);
partial_product_5(333) <= temp_mult_126(333);
partial_product_5(334) <= temp_mult_126(334);
partial_product_5(335) <= temp_mult_126(335);
partial_product_5(336) <= temp_mult_126(336);
partial_product_5(337) <= temp_mult_126(337);
partial_product_5(338) <= temp_mult_132(338);
partial_product_5(339) <= temp_mult_132(339);
partial_product_5(340) <= temp_mult_132(340);
partial_product_5(341) <= temp_mult_132(341);
partial_product_5(342) <= temp_mult_132(342);
partial_product_5(343) <= temp_mult_132(343);
partial_product_5(344) <= temp_mult_132(344);
partial_product_5(345) <= temp_mult_132(345);
partial_product_5(346) <= temp_mult_132(346);
partial_product_5(347) <= temp_mult_132(347);
partial_product_5(348) <= temp_mult_132(348);
partial_product_5(349) <= temp_mult_132(349);
partial_product_5(350) <= temp_mult_132(350);
partial_product_5(351) <= temp_mult_132(351);
partial_product_5(352) <= temp_mult_132(352);
partial_product_5(353) <= temp_mult_132(353);
partial_product_5(354) <= temp_mult_132(354);
partial_product_5(355) <= temp_mult_132(355);
partial_product_5(356) <= temp_mult_132(356);
partial_product_5(357) <= temp_mult_132(357);
partial_product_5(358) <= temp_mult_132(358);
partial_product_5(359) <= temp_mult_132(359);
partial_product_5(360) <= temp_mult_132(360);
partial_product_5(361) <= temp_mult_132(361);
partial_product_5(362) <= temp_mult_132(362);
partial_product_5(363) <= temp_mult_132(363);
partial_product_5(364) <= temp_mult_132(364);
partial_product_5(365) <= temp_mult_132(365);
partial_product_5(366) <= temp_mult_132(366);
partial_product_5(367) <= temp_mult_132(367);
partial_product_5(368) <= temp_mult_132(368);
partial_product_5(369) <= temp_mult_132(369);
partial_product_5(370) <= temp_mult_132(370);
partial_product_5(371) <= temp_mult_132(371);
partial_product_5(372) <= temp_mult_132(372);
partial_product_5(373) <= temp_mult_132(373);
partial_product_5(374) <= temp_mult_132(374);
partial_product_5(375) <= temp_mult_132(375);
partial_product_5(376) <= temp_mult_132(376);
partial_product_5(377) <= temp_mult_132(377);
partial_product_5(378) <= temp_mult_132(378);
partial_product_5(379) <= '0';
partial_product_5(380) <= '0';
partial_product_5(381) <= '0';
partial_product_5(382) <= temp_mult_151(382);
partial_product_5(383) <= temp_mult_151(383);
partial_product_5(384) <= temp_mult_151(384);
partial_product_5(385) <= temp_mult_151(385);
partial_product_5(386) <= temp_mult_151(386);
partial_product_5(387) <= temp_mult_151(387);
partial_product_5(388) <= temp_mult_151(388);
partial_product_5(389) <= temp_mult_151(389);
partial_product_5(390) <= temp_mult_151(390);
partial_product_5(391) <= temp_mult_151(391);
partial_product_5(392) <= temp_mult_151(392);
partial_product_5(393) <= temp_mult_151(393);
partial_product_5(394) <= temp_mult_151(394);
partial_product_5(395) <= temp_mult_151(395);
partial_product_5(396) <= temp_mult_151(396);
partial_product_5(397) <= temp_mult_151(397);
partial_product_5(398) <= temp_mult_151(398);
partial_product_5(399) <= temp_mult_151(399);
partial_product_5(400) <= temp_mult_151(400);
partial_product_5(401) <= temp_mult_151(401);
partial_product_5(402) <= temp_mult_151(402);
partial_product_5(403) <= temp_mult_151(403);
partial_product_5(404) <= temp_mult_151(404);
partial_product_5(405) <= temp_mult_151(405);
partial_product_5(406) <= temp_mult_151(406);
partial_product_5(407) <= temp_mult_151(407);
partial_product_5(408) <= temp_mult_151(408);
partial_product_5(409) <= temp_mult_151(409);
partial_product_5(410) <= temp_mult_151(410);
partial_product_5(411) <= temp_mult_151(411);
partial_product_5(412) <= temp_mult_151(412);
partial_product_5(413) <= temp_mult_151(413);
partial_product_5(414) <= temp_mult_151(414);
partial_product_5(415) <= temp_mult_151(415);
partial_product_5(416) <= temp_mult_151(416);
partial_product_5(417) <= temp_mult_151(417);
partial_product_5(418) <= temp_mult_151(418);
partial_product_5(419) <= temp_mult_151(419);
partial_product_5(420) <= temp_mult_151(420);
partial_product_5(421) <= temp_mult_151(421);
partial_product_5(422) <= temp_mult_151(422);
partial_product_5(423) <= temp_mult_157(423);
partial_product_5(424) <= temp_mult_157(424);
partial_product_5(425) <= temp_mult_157(425);
partial_product_5(426) <= temp_mult_157(426);
partial_product_5(427) <= temp_mult_157(427);
partial_product_5(428) <= temp_mult_157(428);
partial_product_5(429) <= temp_mult_157(429);
partial_product_5(430) <= temp_mult_157(430);
partial_product_5(431) <= temp_mult_157(431);
partial_product_5(432) <= temp_mult_157(432);
partial_product_5(433) <= temp_mult_157(433);
partial_product_5(434) <= temp_mult_157(434);
partial_product_5(435) <= temp_mult_157(435);
partial_product_5(436) <= temp_mult_157(436);
partial_product_5(437) <= temp_mult_157(437);
partial_product_5(438) <= temp_mult_157(438);
partial_product_5(439) <= temp_mult_157(439);
partial_product_5(440) <= temp_mult_157(440);
partial_product_5(441) <= temp_mult_157(441);
partial_product_5(442) <= temp_mult_157(442);
partial_product_5(443) <= temp_mult_157(443);
partial_product_5(444) <= temp_mult_157(444);
partial_product_5(445) <= temp_mult_157(445);
partial_product_5(446) <= temp_mult_157(446);
partial_product_5(447) <= temp_mult_157(447);
partial_product_5(448) <= temp_mult_157(448);
partial_product_5(449) <= temp_mult_157(449);
partial_product_5(450) <= temp_mult_157(450);
partial_product_5(451) <= temp_mult_157(451);
partial_product_5(452) <= temp_mult_157(452);
partial_product_5(453) <= temp_mult_157(453);
partial_product_5(454) <= temp_mult_157(454);
partial_product_5(455) <= temp_mult_157(455);
partial_product_5(456) <= temp_mult_157(456);
partial_product_5(457) <= temp_mult_157(457);
partial_product_5(458) <= temp_mult_157(458);
partial_product_5(459) <= temp_mult_157(459);
partial_product_5(460) <= temp_mult_157(460);
partial_product_5(461) <= temp_mult_157(461);
partial_product_5(462) <= temp_mult_157(462);
partial_product_5(463) <= temp_mult_157(463);
partial_product_5(464) <= '0';
partial_product_5(465) <= '0';
partial_product_5(466) <= '0';
partial_product_5(467) <= '0';
partial_product_5(468) <= '0';
partial_product_5(469) <= '0';
partial_product_5(470) <= '0';
partial_product_5(471) <= '0';
partial_product_5(472) <= '0';
partial_product_5(473) <= '0';
partial_product_5(474) <= '0';
partial_product_5(475) <= '0';
partial_product_5(476) <= '0';
partial_product_5(477) <= '0';
partial_product_5(478) <= '0';
partial_product_5(479) <= '0';
partial_product_5(480) <= '0';
partial_product_5(481) <= '0';
partial_product_5(482) <= '0';
partial_product_5(483) <= '0';
partial_product_5(484) <= '0';
partial_product_5(485) <= '0';
partial_product_5(486) <= '0';
partial_product_5(487) <= '0';
partial_product_5(488) <= '0';
partial_product_5(489) <= '0';
partial_product_5(490) <= '0';
partial_product_5(491) <= '0';
partial_product_5(492) <= '0';
partial_product_5(493) <= '0';
partial_product_5(494) <= '0';
partial_product_5(495) <= '0';
partial_product_5(496) <= '0';
partial_product_5(497) <= '0';
partial_product_5(498) <= '0';
partial_product_5(499) <= '0';
partial_product_5(500) <= '0';
partial_product_5(501) <= '0';
partial_product_5(502) <= '0';
partial_product_5(503) <= '0';
partial_product_5(504) <= '0';
partial_product_5(505) <= '0';
partial_product_5(506) <= '0';
partial_product_5(507) <= '0';
partial_product_5(508) <= '0';
partial_product_5(509) <= '0';
partial_product_5(510) <= '0';
partial_product_5(511) <= '0';
partial_product_5(512) <= '0';
partial_product_6(0) <= '0';
partial_product_6(1) <= '0';
partial_product_6(2) <= '0';
partial_product_6(3) <= '0';
partial_product_6(4) <= '0';
partial_product_6(5) <= '0';
partial_product_6(6) <= '0';
partial_product_6(7) <= '0';
partial_product_6(8) <= '0';
partial_product_6(9) <= '0';
partial_product_6(10) <= '0';
partial_product_6(11) <= '0';
partial_product_6(12) <= '0';
partial_product_6(13) <= '0';
partial_product_6(14) <= '0';
partial_product_6(15) <= '0';
partial_product_6(16) <= '0';
partial_product_6(17) <= '0';
partial_product_6(18) <= '0';
partial_product_6(19) <= '0';
partial_product_6(20) <= '0';
partial_product_6(21) <= '0';
partial_product_6(22) <= '0';
partial_product_6(23) <= '0';
partial_product_6(24) <= '0';
partial_product_6(25) <= '0';
partial_product_6(26) <= '0';
partial_product_6(27) <= '0';
partial_product_6(28) <= '0';
partial_product_6(29) <= '0';
partial_product_6(30) <= '0';
partial_product_6(31) <= '0';
partial_product_6(32) <= '0';
partial_product_6(33) <= '0';
partial_product_6(34) <= '0';
partial_product_6(35) <= '0';
partial_product_6(36) <= '0';
partial_product_6(37) <= '0';
partial_product_6(38) <= '0';
partial_product_6(39) <= '0';
partial_product_6(40) <= '0';
partial_product_6(41) <= '0';
partial_product_6(42) <= '0';
partial_product_6(43) <= '0';
partial_product_6(44) <= '0';
partial_product_6(45) <= '0';
partial_product_6(46) <= '0';
partial_product_6(47) <= '0';
partial_product_6(48) <= '0';
partial_product_6(49) <= '0';
partial_product_6(50) <= '0';
partial_product_6(51) <= '0';
partial_product_6(52) <= '0';
partial_product_6(53) <= '0';
partial_product_6(54) <= '0';
partial_product_6(55) <= '0';
partial_product_6(56) <= '0';
partial_product_6(57) <= '0';
partial_product_6(58) <= '0';
partial_product_6(59) <= '0';
partial_product_6(60) <= '0';
partial_product_6(61) <= '0';
partial_product_6(62) <= '0';
partial_product_6(63) <= '0';
partial_product_6(64) <= '0';
partial_product_6(65) <= '0';
partial_product_6(66) <= '0';
partial_product_6(67) <= '0';
partial_product_6(68) <= temp_mult_20(68);
partial_product_6(69) <= temp_mult_20(69);
partial_product_6(70) <= temp_mult_20(70);
partial_product_6(71) <= temp_mult_20(71);
partial_product_6(72) <= temp_mult_20(72);
partial_product_6(73) <= temp_mult_20(73);
partial_product_6(74) <= temp_mult_20(74);
partial_product_6(75) <= temp_mult_20(75);
partial_product_6(76) <= temp_mult_20(76);
partial_product_6(77) <= temp_mult_20(77);
partial_product_6(78) <= temp_mult_20(78);
partial_product_6(79) <= temp_mult_20(79);
partial_product_6(80) <= temp_mult_20(80);
partial_product_6(81) <= temp_mult_20(81);
partial_product_6(82) <= temp_mult_20(82);
partial_product_6(83) <= temp_mult_20(83);
partial_product_6(84) <= temp_mult_20(84);
partial_product_6(85) <= temp_mult_20(85);
partial_product_6(86) <= temp_mult_20(86);
partial_product_6(87) <= temp_mult_20(87);
partial_product_6(88) <= temp_mult_20(88);
partial_product_6(89) <= temp_mult_20(89);
partial_product_6(90) <= temp_mult_20(90);
partial_product_6(91) <= temp_mult_20(91);
partial_product_6(92) <= temp_mult_20(92);
partial_product_6(93) <= temp_mult_20(93);
partial_product_6(94) <= temp_mult_20(94);
partial_product_6(95) <= temp_mult_20(95);
partial_product_6(96) <= temp_mult_20(96);
partial_product_6(97) <= temp_mult_20(97);
partial_product_6(98) <= temp_mult_20(98);
partial_product_6(99) <= temp_mult_20(99);
partial_product_6(100) <= temp_mult_20(100);
partial_product_6(101) <= temp_mult_20(101);
partial_product_6(102) <= temp_mult_20(102);
partial_product_6(103) <= temp_mult_20(103);
partial_product_6(104) <= temp_mult_20(104);
partial_product_6(105) <= temp_mult_20(105);
partial_product_6(106) <= temp_mult_20(106);
partial_product_6(107) <= temp_mult_20(107);
partial_product_6(108) <= temp_mult_20(108);
partial_product_6(109) <= temp_mult_26(109);
partial_product_6(110) <= temp_mult_26(110);
partial_product_6(111) <= temp_mult_26(111);
partial_product_6(112) <= temp_mult_26(112);
partial_product_6(113) <= temp_mult_26(113);
partial_product_6(114) <= temp_mult_26(114);
partial_product_6(115) <= temp_mult_26(115);
partial_product_6(116) <= temp_mult_26(116);
partial_product_6(117) <= temp_mult_26(117);
partial_product_6(118) <= temp_mult_26(118);
partial_product_6(119) <= temp_mult_26(119);
partial_product_6(120) <= temp_mult_26(120);
partial_product_6(121) <= temp_mult_26(121);
partial_product_6(122) <= temp_mult_26(122);
partial_product_6(123) <= temp_mult_26(123);
partial_product_6(124) <= temp_mult_26(124);
partial_product_6(125) <= temp_mult_26(125);
partial_product_6(126) <= temp_mult_26(126);
partial_product_6(127) <= temp_mult_26(127);
partial_product_6(128) <= temp_mult_26(128);
partial_product_6(129) <= temp_mult_26(129);
partial_product_6(130) <= temp_mult_26(130);
partial_product_6(131) <= temp_mult_26(131);
partial_product_6(132) <= temp_mult_26(132);
partial_product_6(133) <= temp_mult_26(133);
partial_product_6(134) <= temp_mult_26(134);
partial_product_6(135) <= temp_mult_26(135);
partial_product_6(136) <= temp_mult_26(136);
partial_product_6(137) <= temp_mult_26(137);
partial_product_6(138) <= temp_mult_26(138);
partial_product_6(139) <= temp_mult_26(139);
partial_product_6(140) <= temp_mult_26(140);
partial_product_6(141) <= temp_mult_26(141);
partial_product_6(142) <= temp_mult_26(142);
partial_product_6(143) <= temp_mult_26(143);
partial_product_6(144) <= temp_mult_26(144);
partial_product_6(145) <= temp_mult_26(145);
partial_product_6(146) <= temp_mult_26(146);
partial_product_6(147) <= temp_mult_26(147);
partial_product_6(148) <= temp_mult_26(148);
partial_product_6(149) <= temp_mult_26(149);
partial_product_6(150) <= temp_mult_32(150);
partial_product_6(151) <= temp_mult_32(151);
partial_product_6(152) <= temp_mult_32(152);
partial_product_6(153) <= temp_mult_32(153);
partial_product_6(154) <= temp_mult_32(154);
partial_product_6(155) <= temp_mult_32(155);
partial_product_6(156) <= temp_mult_32(156);
partial_product_6(157) <= temp_mult_32(157);
partial_product_6(158) <= temp_mult_32(158);
partial_product_6(159) <= temp_mult_32(159);
partial_product_6(160) <= temp_mult_32(160);
partial_product_6(161) <= temp_mult_32(161);
partial_product_6(162) <= temp_mult_32(162);
partial_product_6(163) <= temp_mult_32(163);
partial_product_6(164) <= temp_mult_32(164);
partial_product_6(165) <= temp_mult_32(165);
partial_product_6(166) <= temp_mult_32(166);
partial_product_6(167) <= temp_mult_32(167);
partial_product_6(168) <= temp_mult_32(168);
partial_product_6(169) <= temp_mult_32(169);
partial_product_6(170) <= temp_mult_32(170);
partial_product_6(171) <= temp_mult_32(171);
partial_product_6(172) <= temp_mult_32(172);
partial_product_6(173) <= temp_mult_32(173);
partial_product_6(174) <= temp_mult_32(174);
partial_product_6(175) <= temp_mult_32(175);
partial_product_6(176) <= temp_mult_32(176);
partial_product_6(177) <= temp_mult_32(177);
partial_product_6(178) <= temp_mult_32(178);
partial_product_6(179) <= temp_mult_32(179);
partial_product_6(180) <= temp_mult_32(180);
partial_product_6(181) <= temp_mult_32(181);
partial_product_6(182) <= temp_mult_32(182);
partial_product_6(183) <= temp_mult_32(183);
partial_product_6(184) <= temp_mult_32(184);
partial_product_6(185) <= temp_mult_32(185);
partial_product_6(186) <= temp_mult_32(186);
partial_product_6(187) <= temp_mult_32(187);
partial_product_6(188) <= temp_mult_32(188);
partial_product_6(189) <= temp_mult_32(189);
partial_product_6(190) <= temp_mult_32(190);
partial_product_6(191) <= temp_mult_38(191);
partial_product_6(192) <= temp_mult_38(192);
partial_product_6(193) <= temp_mult_38(193);
partial_product_6(194) <= temp_mult_38(194);
partial_product_6(195) <= temp_mult_38(195);
partial_product_6(196) <= temp_mult_38(196);
partial_product_6(197) <= temp_mult_38(197);
partial_product_6(198) <= temp_mult_38(198);
partial_product_6(199) <= temp_mult_38(199);
partial_product_6(200) <= temp_mult_38(200);
partial_product_6(201) <= temp_mult_38(201);
partial_product_6(202) <= temp_mult_38(202);
partial_product_6(203) <= temp_mult_38(203);
partial_product_6(204) <= temp_mult_38(204);
partial_product_6(205) <= temp_mult_38(205);
partial_product_6(206) <= temp_mult_38(206);
partial_product_6(207) <= temp_mult_38(207);
partial_product_6(208) <= temp_mult_38(208);
partial_product_6(209) <= temp_mult_38(209);
partial_product_6(210) <= temp_mult_38(210);
partial_product_6(211) <= temp_mult_38(211);
partial_product_6(212) <= temp_mult_38(212);
partial_product_6(213) <= temp_mult_38(213);
partial_product_6(214) <= temp_mult_38(214);
partial_product_6(215) <= temp_mult_38(215);
partial_product_6(216) <= temp_mult_38(216);
partial_product_6(217) <= temp_mult_38(217);
partial_product_6(218) <= temp_mult_38(218);
partial_product_6(219) <= temp_mult_38(219);
partial_product_6(220) <= temp_mult_38(220);
partial_product_6(221) <= temp_mult_38(221);
partial_product_6(222) <= temp_mult_38(222);
partial_product_6(223) <= temp_mult_38(223);
partial_product_6(224) <= temp_mult_38(224);
partial_product_6(225) <= temp_mult_38(225);
partial_product_6(226) <= temp_mult_38(226);
partial_product_6(227) <= temp_mult_38(227);
partial_product_6(228) <= temp_mult_38(228);
partial_product_6(229) <= temp_mult_38(229);
partial_product_6(230) <= temp_mult_38(230);
partial_product_6(231) <= temp_mult_38(231);
partial_product_6(232) <= temp_mult_112(232);
partial_product_6(233) <= temp_mult_112(233);
partial_product_6(234) <= temp_mult_112(234);
partial_product_6(235) <= temp_mult_112(235);
partial_product_6(236) <= temp_mult_112(236);
partial_product_6(237) <= temp_mult_112(237);
partial_product_6(238) <= temp_mult_112(238);
partial_product_6(239) <= temp_mult_112(239);
partial_product_6(240) <= temp_mult_112(240);
partial_product_6(241) <= temp_mult_112(241);
partial_product_6(242) <= temp_mult_112(242);
partial_product_6(243) <= temp_mult_112(243);
partial_product_6(244) <= temp_mult_112(244);
partial_product_6(245) <= temp_mult_112(245);
partial_product_6(246) <= temp_mult_112(246);
partial_product_6(247) <= temp_mult_112(247);
partial_product_6(248) <= temp_mult_112(248);
partial_product_6(249) <= temp_mult_112(249);
partial_product_6(250) <= temp_mult_112(250);
partial_product_6(251) <= temp_mult_112(251);
partial_product_6(252) <= temp_mult_112(252);
partial_product_6(253) <= temp_mult_112(253);
partial_product_6(254) <= temp_mult_112(254);
partial_product_6(255) <= temp_mult_112(255);
partial_product_6(256) <= temp_mult_112(256);
partial_product_6(257) <= temp_mult_112(257);
partial_product_6(258) <= temp_mult_112(258);
partial_product_6(259) <= temp_mult_112(259);
partial_product_6(260) <= temp_mult_112(260);
partial_product_6(261) <= temp_mult_112(261);
partial_product_6(262) <= temp_mult_112(262);
partial_product_6(263) <= temp_mult_112(263);
partial_product_6(264) <= temp_mult_112(264);
partial_product_6(265) <= temp_mult_112(265);
partial_product_6(266) <= temp_mult_112(266);
partial_product_6(267) <= temp_mult_112(267);
partial_product_6(268) <= temp_mult_112(268);
partial_product_6(269) <= temp_mult_112(269);
partial_product_6(270) <= temp_mult_112(270);
partial_product_6(271) <= temp_mult_112(271);
partial_product_6(272) <= temp_mult_112(272);
partial_product_6(273) <= temp_mult_125(273);
partial_product_6(274) <= temp_mult_125(274);
partial_product_6(275) <= temp_mult_125(275);
partial_product_6(276) <= temp_mult_125(276);
partial_product_6(277) <= temp_mult_125(277);
partial_product_6(278) <= temp_mult_125(278);
partial_product_6(279) <= temp_mult_125(279);
partial_product_6(280) <= temp_mult_125(280);
partial_product_6(281) <= temp_mult_125(281);
partial_product_6(282) <= temp_mult_125(282);
partial_product_6(283) <= temp_mult_125(283);
partial_product_6(284) <= temp_mult_125(284);
partial_product_6(285) <= temp_mult_125(285);
partial_product_6(286) <= temp_mult_125(286);
partial_product_6(287) <= temp_mult_125(287);
partial_product_6(288) <= temp_mult_125(288);
partial_product_6(289) <= temp_mult_125(289);
partial_product_6(290) <= temp_mult_125(290);
partial_product_6(291) <= temp_mult_125(291);
partial_product_6(292) <= temp_mult_125(292);
partial_product_6(293) <= temp_mult_125(293);
partial_product_6(294) <= temp_mult_125(294);
partial_product_6(295) <= temp_mult_125(295);
partial_product_6(296) <= temp_mult_125(296);
partial_product_6(297) <= temp_mult_125(297);
partial_product_6(298) <= temp_mult_125(298);
partial_product_6(299) <= temp_mult_125(299);
partial_product_6(300) <= temp_mult_125(300);
partial_product_6(301) <= temp_mult_125(301);
partial_product_6(302) <= temp_mult_125(302);
partial_product_6(303) <= temp_mult_125(303);
partial_product_6(304) <= temp_mult_125(304);
partial_product_6(305) <= temp_mult_125(305);
partial_product_6(306) <= temp_mult_125(306);
partial_product_6(307) <= temp_mult_125(307);
partial_product_6(308) <= temp_mult_125(308);
partial_product_6(309) <= temp_mult_125(309);
partial_product_6(310) <= temp_mult_125(310);
partial_product_6(311) <= temp_mult_125(311);
partial_product_6(312) <= temp_mult_125(312);
partial_product_6(313) <= temp_mult_125(313);
partial_product_6(314) <= temp_mult_131(314);
partial_product_6(315) <= temp_mult_131(315);
partial_product_6(316) <= temp_mult_131(316);
partial_product_6(317) <= temp_mult_131(317);
partial_product_6(318) <= temp_mult_131(318);
partial_product_6(319) <= temp_mult_131(319);
partial_product_6(320) <= temp_mult_131(320);
partial_product_6(321) <= temp_mult_131(321);
partial_product_6(322) <= temp_mult_131(322);
partial_product_6(323) <= temp_mult_131(323);
partial_product_6(324) <= temp_mult_131(324);
partial_product_6(325) <= temp_mult_131(325);
partial_product_6(326) <= temp_mult_131(326);
partial_product_6(327) <= temp_mult_131(327);
partial_product_6(328) <= temp_mult_131(328);
partial_product_6(329) <= temp_mult_131(329);
partial_product_6(330) <= temp_mult_131(330);
partial_product_6(331) <= temp_mult_131(331);
partial_product_6(332) <= temp_mult_131(332);
partial_product_6(333) <= temp_mult_131(333);
partial_product_6(334) <= temp_mult_131(334);
partial_product_6(335) <= temp_mult_131(335);
partial_product_6(336) <= temp_mult_131(336);
partial_product_6(337) <= temp_mult_131(337);
partial_product_6(338) <= temp_mult_131(338);
partial_product_6(339) <= temp_mult_131(339);
partial_product_6(340) <= temp_mult_131(340);
partial_product_6(341) <= temp_mult_131(341);
partial_product_6(342) <= temp_mult_131(342);
partial_product_6(343) <= temp_mult_131(343);
partial_product_6(344) <= temp_mult_131(344);
partial_product_6(345) <= temp_mult_131(345);
partial_product_6(346) <= temp_mult_131(346);
partial_product_6(347) <= temp_mult_131(347);
partial_product_6(348) <= temp_mult_131(348);
partial_product_6(349) <= temp_mult_131(349);
partial_product_6(350) <= temp_mult_131(350);
partial_product_6(351) <= temp_mult_131(351);
partial_product_6(352) <= temp_mult_131(352);
partial_product_6(353) <= temp_mult_131(353);
partial_product_6(354) <= temp_mult_131(354);
partial_product_6(355) <= temp_mult_137(355);
partial_product_6(356) <= temp_mult_137(356);
partial_product_6(357) <= temp_mult_137(357);
partial_product_6(358) <= temp_mult_137(358);
partial_product_6(359) <= temp_mult_137(359);
partial_product_6(360) <= temp_mult_137(360);
partial_product_6(361) <= temp_mult_137(361);
partial_product_6(362) <= temp_mult_137(362);
partial_product_6(363) <= temp_mult_137(363);
partial_product_6(364) <= temp_mult_137(364);
partial_product_6(365) <= temp_mult_137(365);
partial_product_6(366) <= temp_mult_137(366);
partial_product_6(367) <= temp_mult_137(367);
partial_product_6(368) <= temp_mult_137(368);
partial_product_6(369) <= temp_mult_137(369);
partial_product_6(370) <= temp_mult_137(370);
partial_product_6(371) <= temp_mult_137(371);
partial_product_6(372) <= temp_mult_137(372);
partial_product_6(373) <= temp_mult_137(373);
partial_product_6(374) <= temp_mult_137(374);
partial_product_6(375) <= temp_mult_137(375);
partial_product_6(376) <= temp_mult_137(376);
partial_product_6(377) <= temp_mult_137(377);
partial_product_6(378) <= temp_mult_137(378);
partial_product_6(379) <= temp_mult_137(379);
partial_product_6(380) <= temp_mult_137(380);
partial_product_6(381) <= temp_mult_137(381);
partial_product_6(382) <= temp_mult_137(382);
partial_product_6(383) <= temp_mult_137(383);
partial_product_6(384) <= temp_mult_137(384);
partial_product_6(385) <= temp_mult_137(385);
partial_product_6(386) <= temp_mult_137(386);
partial_product_6(387) <= temp_mult_137(387);
partial_product_6(388) <= temp_mult_137(388);
partial_product_6(389) <= temp_mult_137(389);
partial_product_6(390) <= temp_mult_137(390);
partial_product_6(391) <= temp_mult_137(391);
partial_product_6(392) <= temp_mult_137(392);
partial_product_6(393) <= temp_mult_137(393);
partial_product_6(394) <= temp_mult_137(394);
partial_product_6(395) <= temp_mult_137(395);
partial_product_6(396) <= '0';
partial_product_6(397) <= '0';
partial_product_6(398) <= '0';
partial_product_6(399) <= temp_mult_156(399);
partial_product_6(400) <= temp_mult_156(400);
partial_product_6(401) <= temp_mult_156(401);
partial_product_6(402) <= temp_mult_156(402);
partial_product_6(403) <= temp_mult_156(403);
partial_product_6(404) <= temp_mult_156(404);
partial_product_6(405) <= temp_mult_156(405);
partial_product_6(406) <= temp_mult_156(406);
partial_product_6(407) <= temp_mult_156(407);
partial_product_6(408) <= temp_mult_156(408);
partial_product_6(409) <= temp_mult_156(409);
partial_product_6(410) <= temp_mult_156(410);
partial_product_6(411) <= temp_mult_156(411);
partial_product_6(412) <= temp_mult_156(412);
partial_product_6(413) <= temp_mult_156(413);
partial_product_6(414) <= temp_mult_156(414);
partial_product_6(415) <= temp_mult_156(415);
partial_product_6(416) <= temp_mult_156(416);
partial_product_6(417) <= temp_mult_156(417);
partial_product_6(418) <= temp_mult_156(418);
partial_product_6(419) <= temp_mult_156(419);
partial_product_6(420) <= temp_mult_156(420);
partial_product_6(421) <= temp_mult_156(421);
partial_product_6(422) <= temp_mult_156(422);
partial_product_6(423) <= temp_mult_156(423);
partial_product_6(424) <= temp_mult_156(424);
partial_product_6(425) <= temp_mult_156(425);
partial_product_6(426) <= temp_mult_156(426);
partial_product_6(427) <= temp_mult_156(427);
partial_product_6(428) <= temp_mult_156(428);
partial_product_6(429) <= temp_mult_156(429);
partial_product_6(430) <= temp_mult_156(430);
partial_product_6(431) <= temp_mult_156(431);
partial_product_6(432) <= temp_mult_156(432);
partial_product_6(433) <= temp_mult_156(433);
partial_product_6(434) <= temp_mult_156(434);
partial_product_6(435) <= temp_mult_156(435);
partial_product_6(436) <= temp_mult_156(436);
partial_product_6(437) <= temp_mult_156(437);
partial_product_6(438) <= temp_mult_156(438);
partial_product_6(439) <= temp_mult_156(439);
partial_product_6(440) <= '0';
partial_product_6(441) <= '0';
partial_product_6(442) <= '0';
partial_product_6(443) <= '0';
partial_product_6(444) <= '0';
partial_product_6(445) <= '0';
partial_product_6(446) <= '0';
partial_product_6(447) <= '0';
partial_product_6(448) <= '0';
partial_product_6(449) <= '0';
partial_product_6(450) <= '0';
partial_product_6(451) <= '0';
partial_product_6(452) <= '0';
partial_product_6(453) <= '0';
partial_product_6(454) <= '0';
partial_product_6(455) <= '0';
partial_product_6(456) <= '0';
partial_product_6(457) <= '0';
partial_product_6(458) <= '0';
partial_product_6(459) <= '0';
partial_product_6(460) <= '0';
partial_product_6(461) <= '0';
partial_product_6(462) <= '0';
partial_product_6(463) <= '0';
partial_product_6(464) <= '0';
partial_product_6(465) <= '0';
partial_product_6(466) <= '0';
partial_product_6(467) <= '0';
partial_product_6(468) <= '0';
partial_product_6(469) <= '0';
partial_product_6(470) <= '0';
partial_product_6(471) <= '0';
partial_product_6(472) <= '0';
partial_product_6(473) <= '0';
partial_product_6(474) <= '0';
partial_product_6(475) <= '0';
partial_product_6(476) <= '0';
partial_product_6(477) <= '0';
partial_product_6(478) <= '0';
partial_product_6(479) <= '0';
partial_product_6(480) <= '0';
partial_product_6(481) <= '0';
partial_product_6(482) <= '0';
partial_product_6(483) <= '0';
partial_product_6(484) <= '0';
partial_product_6(485) <= '0';
partial_product_6(486) <= '0';
partial_product_6(487) <= '0';
partial_product_6(488) <= '0';
partial_product_6(489) <= '0';
partial_product_6(490) <= '0';
partial_product_6(491) <= '0';
partial_product_6(492) <= '0';
partial_product_6(493) <= '0';
partial_product_6(494) <= '0';
partial_product_6(495) <= '0';
partial_product_6(496) <= '0';
partial_product_6(497) <= '0';
partial_product_6(498) <= '0';
partial_product_6(499) <= '0';
partial_product_6(500) <= '0';
partial_product_6(501) <= '0';
partial_product_6(502) <= '0';
partial_product_6(503) <= '0';
partial_product_6(504) <= '0';
partial_product_6(505) <= '0';
partial_product_6(506) <= '0';
partial_product_6(507) <= '0';
partial_product_6(508) <= '0';
partial_product_6(509) <= '0';
partial_product_6(510) <= '0';
partial_product_6(511) <= '0';
partial_product_6(512) <= '0';
partial_product_7(0) <= '0';
partial_product_7(1) <= '0';
partial_product_7(2) <= '0';
partial_product_7(3) <= '0';
partial_product_7(4) <= '0';
partial_product_7(5) <= '0';
partial_product_7(6) <= '0';
partial_product_7(7) <= '0';
partial_product_7(8) <= '0';
partial_product_7(9) <= '0';
partial_product_7(10) <= '0';
partial_product_7(11) <= '0';
partial_product_7(12) <= '0';
partial_product_7(13) <= '0';
partial_product_7(14) <= '0';
partial_product_7(15) <= '0';
partial_product_7(16) <= '0';
partial_product_7(17) <= '0';
partial_product_7(18) <= '0';
partial_product_7(19) <= '0';
partial_product_7(20) <= '0';
partial_product_7(21) <= '0';
partial_product_7(22) <= '0';
partial_product_7(23) <= '0';
partial_product_7(24) <= '0';
partial_product_7(25) <= '0';
partial_product_7(26) <= '0';
partial_product_7(27) <= '0';
partial_product_7(28) <= '0';
partial_product_7(29) <= '0';
partial_product_7(30) <= '0';
partial_product_7(31) <= '0';
partial_product_7(32) <= '0';
partial_product_7(33) <= '0';
partial_product_7(34) <= '0';
partial_product_7(35) <= '0';
partial_product_7(36) <= '0';
partial_product_7(37) <= '0';
partial_product_7(38) <= '0';
partial_product_7(39) <= '0';
partial_product_7(40) <= '0';
partial_product_7(41) <= '0';
partial_product_7(42) <= '0';
partial_product_7(43) <= '0';
partial_product_7(44) <= '0';
partial_product_7(45) <= '0';
partial_product_7(46) <= '0';
partial_product_7(47) <= '0';
partial_product_7(48) <= '0';
partial_product_7(49) <= '0';
partial_product_7(50) <= '0';
partial_product_7(51) <= '0';
partial_product_7(52) <= '0';
partial_product_7(53) <= '0';
partial_product_7(54) <= '0';
partial_product_7(55) <= '0';
partial_product_7(56) <= '0';
partial_product_7(57) <= '0';
partial_product_7(58) <= '0';
partial_product_7(59) <= '0';
partial_product_7(60) <= '0';
partial_product_7(61) <= '0';
partial_product_7(62) <= '0';
partial_product_7(63) <= '0';
partial_product_7(64) <= '0';
partial_product_7(65) <= '0';
partial_product_7(66) <= '0';
partial_product_7(67) <= '0';
partial_product_7(68) <= '0';
partial_product_7(69) <= '0';
partial_product_7(70) <= '0';
partial_product_7(71) <= '0';
partial_product_7(72) <= temp_mult_3(72);
partial_product_7(73) <= temp_mult_3(73);
partial_product_7(74) <= temp_mult_3(74);
partial_product_7(75) <= temp_mult_3(75);
partial_product_7(76) <= temp_mult_3(76);
partial_product_7(77) <= temp_mult_3(77);
partial_product_7(78) <= temp_mult_3(78);
partial_product_7(79) <= temp_mult_3(79);
partial_product_7(80) <= temp_mult_3(80);
partial_product_7(81) <= temp_mult_3(81);
partial_product_7(82) <= temp_mult_3(82);
partial_product_7(83) <= temp_mult_3(83);
partial_product_7(84) <= temp_mult_3(84);
partial_product_7(85) <= temp_mult_3(85);
partial_product_7(86) <= temp_mult_3(86);
partial_product_7(87) <= temp_mult_3(87);
partial_product_7(88) <= temp_mult_3(88);
partial_product_7(89) <= temp_mult_3(89);
partial_product_7(90) <= temp_mult_3(90);
partial_product_7(91) <= temp_mult_3(91);
partial_product_7(92) <= temp_mult_3(92);
partial_product_7(93) <= temp_mult_3(93);
partial_product_7(94) <= temp_mult_3(94);
partial_product_7(95) <= temp_mult_3(95);
partial_product_7(96) <= temp_mult_3(96);
partial_product_7(97) <= temp_mult_3(97);
partial_product_7(98) <= temp_mult_3(98);
partial_product_7(99) <= temp_mult_3(99);
partial_product_7(100) <= temp_mult_3(100);
partial_product_7(101) <= temp_mult_3(101);
partial_product_7(102) <= temp_mult_3(102);
partial_product_7(103) <= temp_mult_3(103);
partial_product_7(104) <= temp_mult_3(104);
partial_product_7(105) <= temp_mult_3(105);
partial_product_7(106) <= temp_mult_3(106);
partial_product_7(107) <= temp_mult_3(107);
partial_product_7(108) <= temp_mult_3(108);
partial_product_7(109) <= temp_mult_3(109);
partial_product_7(110) <= temp_mult_3(110);
partial_product_7(111) <= temp_mult_3(111);
partial_product_7(112) <= temp_mult_3(112);
partial_product_7(113) <= temp_mult_9(113);
partial_product_7(114) <= temp_mult_9(114);
partial_product_7(115) <= temp_mult_9(115);
partial_product_7(116) <= temp_mult_9(116);
partial_product_7(117) <= temp_mult_9(117);
partial_product_7(118) <= temp_mult_9(118);
partial_product_7(119) <= temp_mult_9(119);
partial_product_7(120) <= temp_mult_9(120);
partial_product_7(121) <= temp_mult_9(121);
partial_product_7(122) <= temp_mult_9(122);
partial_product_7(123) <= temp_mult_9(123);
partial_product_7(124) <= temp_mult_9(124);
partial_product_7(125) <= temp_mult_9(125);
partial_product_7(126) <= temp_mult_9(126);
partial_product_7(127) <= temp_mult_9(127);
partial_product_7(128) <= temp_mult_9(128);
partial_product_7(129) <= temp_mult_9(129);
partial_product_7(130) <= temp_mult_9(130);
partial_product_7(131) <= temp_mult_9(131);
partial_product_7(132) <= temp_mult_9(132);
partial_product_7(133) <= temp_mult_9(133);
partial_product_7(134) <= temp_mult_9(134);
partial_product_7(135) <= temp_mult_9(135);
partial_product_7(136) <= temp_mult_9(136);
partial_product_7(137) <= temp_mult_9(137);
partial_product_7(138) <= temp_mult_9(138);
partial_product_7(139) <= temp_mult_9(139);
partial_product_7(140) <= temp_mult_9(140);
partial_product_7(141) <= temp_mult_9(141);
partial_product_7(142) <= temp_mult_9(142);
partial_product_7(143) <= temp_mult_9(143);
partial_product_7(144) <= temp_mult_9(144);
partial_product_7(145) <= temp_mult_9(145);
partial_product_7(146) <= temp_mult_9(146);
partial_product_7(147) <= temp_mult_9(147);
partial_product_7(148) <= temp_mult_9(148);
partial_product_7(149) <= temp_mult_9(149);
partial_product_7(150) <= temp_mult_9(150);
partial_product_7(151) <= temp_mult_9(151);
partial_product_7(152) <= temp_mult_9(152);
partial_product_7(153) <= temp_mult_9(153);
partial_product_7(154) <= temp_mult_42(154);
partial_product_7(155) <= temp_mult_42(155);
partial_product_7(156) <= temp_mult_42(156);
partial_product_7(157) <= temp_mult_42(157);
partial_product_7(158) <= temp_mult_42(158);
partial_product_7(159) <= temp_mult_42(159);
partial_product_7(160) <= temp_mult_42(160);
partial_product_7(161) <= temp_mult_42(161);
partial_product_7(162) <= temp_mult_42(162);
partial_product_7(163) <= temp_mult_42(163);
partial_product_7(164) <= temp_mult_42(164);
partial_product_7(165) <= temp_mult_42(165);
partial_product_7(166) <= temp_mult_42(166);
partial_product_7(167) <= temp_mult_42(167);
partial_product_7(168) <= temp_mult_42(168);
partial_product_7(169) <= temp_mult_42(169);
partial_product_7(170) <= temp_mult_42(170);
partial_product_7(171) <= temp_mult_42(171);
partial_product_7(172) <= temp_mult_42(172);
partial_product_7(173) <= temp_mult_42(173);
partial_product_7(174) <= temp_mult_42(174);
partial_product_7(175) <= temp_mult_42(175);
partial_product_7(176) <= temp_mult_42(176);
partial_product_7(177) <= temp_mult_42(177);
partial_product_7(178) <= temp_mult_42(178);
partial_product_7(179) <= temp_mult_42(179);
partial_product_7(180) <= temp_mult_42(180);
partial_product_7(181) <= temp_mult_42(181);
partial_product_7(182) <= temp_mult_42(182);
partial_product_7(183) <= temp_mult_42(183);
partial_product_7(184) <= temp_mult_42(184);
partial_product_7(185) <= temp_mult_42(185);
partial_product_7(186) <= temp_mult_42(186);
partial_product_7(187) <= temp_mult_42(187);
partial_product_7(188) <= temp_mult_42(188);
partial_product_7(189) <= temp_mult_42(189);
partial_product_7(190) <= temp_mult_42(190);
partial_product_7(191) <= temp_mult_42(191);
partial_product_7(192) <= temp_mult_42(192);
partial_product_7(193) <= temp_mult_42(193);
partial_product_7(194) <= temp_mult_42(194);
partial_product_7(195) <= temp_mult_51(195);
partial_product_7(196) <= temp_mult_51(196);
partial_product_7(197) <= temp_mult_51(197);
partial_product_7(198) <= temp_mult_51(198);
partial_product_7(199) <= temp_mult_51(199);
partial_product_7(200) <= temp_mult_51(200);
partial_product_7(201) <= temp_mult_51(201);
partial_product_7(202) <= temp_mult_51(202);
partial_product_7(203) <= temp_mult_51(203);
partial_product_7(204) <= temp_mult_51(204);
partial_product_7(205) <= temp_mult_51(205);
partial_product_7(206) <= temp_mult_51(206);
partial_product_7(207) <= temp_mult_51(207);
partial_product_7(208) <= temp_mult_51(208);
partial_product_7(209) <= temp_mult_51(209);
partial_product_7(210) <= temp_mult_51(210);
partial_product_7(211) <= temp_mult_51(211);
partial_product_7(212) <= temp_mult_51(212);
partial_product_7(213) <= temp_mult_51(213);
partial_product_7(214) <= temp_mult_51(214);
partial_product_7(215) <= temp_mult_51(215);
partial_product_7(216) <= temp_mult_51(216);
partial_product_7(217) <= temp_mult_51(217);
partial_product_7(218) <= temp_mult_51(218);
partial_product_7(219) <= temp_mult_51(219);
partial_product_7(220) <= temp_mult_51(220);
partial_product_7(221) <= temp_mult_51(221);
partial_product_7(222) <= temp_mult_51(222);
partial_product_7(223) <= temp_mult_51(223);
partial_product_7(224) <= temp_mult_51(224);
partial_product_7(225) <= temp_mult_51(225);
partial_product_7(226) <= temp_mult_51(226);
partial_product_7(227) <= temp_mult_51(227);
partial_product_7(228) <= temp_mult_51(228);
partial_product_7(229) <= temp_mult_51(229);
partial_product_7(230) <= temp_mult_51(230);
partial_product_7(231) <= temp_mult_51(231);
partial_product_7(232) <= temp_mult_51(232);
partial_product_7(233) <= temp_mult_51(233);
partial_product_7(234) <= temp_mult_51(234);
partial_product_7(235) <= temp_mult_51(235);
partial_product_7(236) <= temp_mult_60(236);
partial_product_7(237) <= temp_mult_60(237);
partial_product_7(238) <= temp_mult_60(238);
partial_product_7(239) <= temp_mult_60(239);
partial_product_7(240) <= temp_mult_60(240);
partial_product_7(241) <= temp_mult_60(241);
partial_product_7(242) <= temp_mult_60(242);
partial_product_7(243) <= temp_mult_60(243);
partial_product_7(244) <= temp_mult_60(244);
partial_product_7(245) <= temp_mult_60(245);
partial_product_7(246) <= temp_mult_60(246);
partial_product_7(247) <= temp_mult_60(247);
partial_product_7(248) <= temp_mult_60(248);
partial_product_7(249) <= temp_mult_60(249);
partial_product_7(250) <= temp_mult_60(250);
partial_product_7(251) <= temp_mult_60(251);
partial_product_7(252) <= temp_mult_60(252);
partial_product_7(253) <= temp_mult_60(253);
partial_product_7(254) <= temp_mult_60(254);
partial_product_7(255) <= temp_mult_60(255);
partial_product_7(256) <= temp_mult_60(256);
partial_product_7(257) <= temp_mult_60(257);
partial_product_7(258) <= temp_mult_60(258);
partial_product_7(259) <= temp_mult_60(259);
partial_product_7(260) <= temp_mult_60(260);
partial_product_7(261) <= temp_mult_60(261);
partial_product_7(262) <= temp_mult_60(262);
partial_product_7(263) <= temp_mult_60(263);
partial_product_7(264) <= temp_mult_60(264);
partial_product_7(265) <= temp_mult_60(265);
partial_product_7(266) <= temp_mult_60(266);
partial_product_7(267) <= temp_mult_60(267);
partial_product_7(268) <= temp_mult_60(268);
partial_product_7(269) <= temp_mult_60(269);
partial_product_7(270) <= temp_mult_60(270);
partial_product_7(271) <= temp_mult_60(271);
partial_product_7(272) <= temp_mult_60(272);
partial_product_7(273) <= temp_mult_60(273);
partial_product_7(274) <= temp_mult_60(274);
partial_product_7(275) <= temp_mult_60(275);
partial_product_7(276) <= temp_mult_60(276);
partial_product_7(277) <= temp_mult_69(277);
partial_product_7(278) <= temp_mult_69(278);
partial_product_7(279) <= temp_mult_69(279);
partial_product_7(280) <= temp_mult_69(280);
partial_product_7(281) <= temp_mult_69(281);
partial_product_7(282) <= temp_mult_69(282);
partial_product_7(283) <= temp_mult_69(283);
partial_product_7(284) <= temp_mult_69(284);
partial_product_7(285) <= temp_mult_69(285);
partial_product_7(286) <= temp_mult_69(286);
partial_product_7(287) <= temp_mult_69(287);
partial_product_7(288) <= temp_mult_69(288);
partial_product_7(289) <= temp_mult_69(289);
partial_product_7(290) <= temp_mult_69(290);
partial_product_7(291) <= temp_mult_69(291);
partial_product_7(292) <= temp_mult_69(292);
partial_product_7(293) <= temp_mult_69(293);
partial_product_7(294) <= temp_mult_69(294);
partial_product_7(295) <= temp_mult_69(295);
partial_product_7(296) <= temp_mult_69(296);
partial_product_7(297) <= temp_mult_69(297);
partial_product_7(298) <= temp_mult_69(298);
partial_product_7(299) <= temp_mult_69(299);
partial_product_7(300) <= temp_mult_69(300);
partial_product_7(301) <= temp_mult_69(301);
partial_product_7(302) <= temp_mult_69(302);
partial_product_7(303) <= temp_mult_69(303);
partial_product_7(304) <= temp_mult_69(304);
partial_product_7(305) <= temp_mult_69(305);
partial_product_7(306) <= temp_mult_69(306);
partial_product_7(307) <= temp_mult_69(307);
partial_product_7(308) <= temp_mult_69(308);
partial_product_7(309) <= temp_mult_69(309);
partial_product_7(310) <= temp_mult_69(310);
partial_product_7(311) <= temp_mult_69(311);
partial_product_7(312) <= temp_mult_69(312);
partial_product_7(313) <= temp_mult_69(313);
partial_product_7(314) <= temp_mult_69(314);
partial_product_7(315) <= temp_mult_69(315);
partial_product_7(316) <= temp_mult_69(316);
partial_product_7(317) <= temp_mult_69(317);
partial_product_7(318) <= temp_mult_78(318);
partial_product_7(319) <= temp_mult_78(319);
partial_product_7(320) <= temp_mult_78(320);
partial_product_7(321) <= temp_mult_78(321);
partial_product_7(322) <= temp_mult_78(322);
partial_product_7(323) <= temp_mult_78(323);
partial_product_7(324) <= temp_mult_78(324);
partial_product_7(325) <= temp_mult_78(325);
partial_product_7(326) <= temp_mult_78(326);
partial_product_7(327) <= temp_mult_78(327);
partial_product_7(328) <= temp_mult_78(328);
partial_product_7(329) <= temp_mult_78(329);
partial_product_7(330) <= temp_mult_78(330);
partial_product_7(331) <= temp_mult_78(331);
partial_product_7(332) <= temp_mult_78(332);
partial_product_7(333) <= temp_mult_78(333);
partial_product_7(334) <= temp_mult_78(334);
partial_product_7(335) <= temp_mult_78(335);
partial_product_7(336) <= temp_mult_78(336);
partial_product_7(337) <= temp_mult_78(337);
partial_product_7(338) <= temp_mult_78(338);
partial_product_7(339) <= temp_mult_78(339);
partial_product_7(340) <= temp_mult_78(340);
partial_product_7(341) <= temp_mult_78(341);
partial_product_7(342) <= temp_mult_78(342);
partial_product_7(343) <= temp_mult_78(343);
partial_product_7(344) <= temp_mult_78(344);
partial_product_7(345) <= temp_mult_78(345);
partial_product_7(346) <= temp_mult_78(346);
partial_product_7(347) <= temp_mult_78(347);
partial_product_7(348) <= temp_mult_78(348);
partial_product_7(349) <= temp_mult_78(349);
partial_product_7(350) <= temp_mult_78(350);
partial_product_7(351) <= temp_mult_78(351);
partial_product_7(352) <= temp_mult_78(352);
partial_product_7(353) <= temp_mult_78(353);
partial_product_7(354) <= temp_mult_78(354);
partial_product_7(355) <= temp_mult_78(355);
partial_product_7(356) <= temp_mult_78(356);
partial_product_7(357) <= temp_mult_78(357);
partial_product_7(358) <= temp_mult_78(358);
partial_product_7(359) <= '0';
partial_product_7(360) <= '0';
partial_product_7(361) <= '0';
partial_product_7(362) <= '0';
partial_product_7(363) <= '0';
partial_product_7(364) <= '0';
partial_product_7(365) <= temp_mult_146(365);
partial_product_7(366) <= temp_mult_146(366);
partial_product_7(367) <= temp_mult_146(367);
partial_product_7(368) <= temp_mult_146(368);
partial_product_7(369) <= temp_mult_146(369);
partial_product_7(370) <= temp_mult_146(370);
partial_product_7(371) <= temp_mult_146(371);
partial_product_7(372) <= temp_mult_146(372);
partial_product_7(373) <= temp_mult_146(373);
partial_product_7(374) <= temp_mult_146(374);
partial_product_7(375) <= temp_mult_146(375);
partial_product_7(376) <= temp_mult_146(376);
partial_product_7(377) <= temp_mult_146(377);
partial_product_7(378) <= temp_mult_146(378);
partial_product_7(379) <= temp_mult_146(379);
partial_product_7(380) <= temp_mult_146(380);
partial_product_7(381) <= temp_mult_146(381);
partial_product_7(382) <= temp_mult_146(382);
partial_product_7(383) <= temp_mult_146(383);
partial_product_7(384) <= temp_mult_146(384);
partial_product_7(385) <= temp_mult_146(385);
partial_product_7(386) <= temp_mult_146(386);
partial_product_7(387) <= temp_mult_146(387);
partial_product_7(388) <= temp_mult_146(388);
partial_product_7(389) <= temp_mult_146(389);
partial_product_7(390) <= temp_mult_146(390);
partial_product_7(391) <= temp_mult_146(391);
partial_product_7(392) <= temp_mult_146(392);
partial_product_7(393) <= temp_mult_146(393);
partial_product_7(394) <= temp_mult_146(394);
partial_product_7(395) <= temp_mult_146(395);
partial_product_7(396) <= temp_mult_146(396);
partial_product_7(397) <= temp_mult_146(397);
partial_product_7(398) <= temp_mult_146(398);
partial_product_7(399) <= temp_mult_146(399);
partial_product_7(400) <= temp_mult_146(400);
partial_product_7(401) <= temp_mult_146(401);
partial_product_7(402) <= temp_mult_146(402);
partial_product_7(403) <= temp_mult_146(403);
partial_product_7(404) <= temp_mult_146(404);
partial_product_7(405) <= temp_mult_146(405);
partial_product_7(406) <= temp_mult_152(406);
partial_product_7(407) <= temp_mult_152(407);
partial_product_7(408) <= temp_mult_152(408);
partial_product_7(409) <= temp_mult_152(409);
partial_product_7(410) <= temp_mult_152(410);
partial_product_7(411) <= temp_mult_152(411);
partial_product_7(412) <= temp_mult_152(412);
partial_product_7(413) <= temp_mult_152(413);
partial_product_7(414) <= temp_mult_152(414);
partial_product_7(415) <= temp_mult_152(415);
partial_product_7(416) <= temp_mult_152(416);
partial_product_7(417) <= temp_mult_152(417);
partial_product_7(418) <= temp_mult_152(418);
partial_product_7(419) <= temp_mult_152(419);
partial_product_7(420) <= temp_mult_152(420);
partial_product_7(421) <= temp_mult_152(421);
partial_product_7(422) <= temp_mult_152(422);
partial_product_7(423) <= temp_mult_152(423);
partial_product_7(424) <= temp_mult_152(424);
partial_product_7(425) <= temp_mult_152(425);
partial_product_7(426) <= temp_mult_152(426);
partial_product_7(427) <= temp_mult_152(427);
partial_product_7(428) <= temp_mult_152(428);
partial_product_7(429) <= temp_mult_152(429);
partial_product_7(430) <= temp_mult_152(430);
partial_product_7(431) <= temp_mult_152(431);
partial_product_7(432) <= temp_mult_152(432);
partial_product_7(433) <= temp_mult_152(433);
partial_product_7(434) <= temp_mult_152(434);
partial_product_7(435) <= temp_mult_152(435);
partial_product_7(436) <= temp_mult_152(436);
partial_product_7(437) <= temp_mult_152(437);
partial_product_7(438) <= temp_mult_152(438);
partial_product_7(439) <= temp_mult_152(439);
partial_product_7(440) <= temp_mult_152(440);
partial_product_7(441) <= temp_mult_152(441);
partial_product_7(442) <= temp_mult_152(442);
partial_product_7(443) <= temp_mult_152(443);
partial_product_7(444) <= temp_mult_152(444);
partial_product_7(445) <= temp_mult_152(445);
partial_product_7(446) <= temp_mult_152(446);
partial_product_7(447) <= '0';
partial_product_7(448) <= '0';
partial_product_7(449) <= '0';
partial_product_7(450) <= '0';
partial_product_7(451) <= '0';
partial_product_7(452) <= '0';
partial_product_7(453) <= '0';
partial_product_7(454) <= '0';
partial_product_7(455) <= '0';
partial_product_7(456) <= '0';
partial_product_7(457) <= '0';
partial_product_7(458) <= '0';
partial_product_7(459) <= '0';
partial_product_7(460) <= '0';
partial_product_7(461) <= '0';
partial_product_7(462) <= '0';
partial_product_7(463) <= '0';
partial_product_7(464) <= '0';
partial_product_7(465) <= '0';
partial_product_7(466) <= '0';
partial_product_7(467) <= '0';
partial_product_7(468) <= '0';
partial_product_7(469) <= '0';
partial_product_7(470) <= '0';
partial_product_7(471) <= '0';
partial_product_7(472) <= '0';
partial_product_7(473) <= '0';
partial_product_7(474) <= '0';
partial_product_7(475) <= '0';
partial_product_7(476) <= '0';
partial_product_7(477) <= '0';
partial_product_7(478) <= '0';
partial_product_7(479) <= '0';
partial_product_7(480) <= '0';
partial_product_7(481) <= '0';
partial_product_7(482) <= '0';
partial_product_7(483) <= '0';
partial_product_7(484) <= '0';
partial_product_7(485) <= '0';
partial_product_7(486) <= '0';
partial_product_7(487) <= '0';
partial_product_7(488) <= '0';
partial_product_7(489) <= '0';
partial_product_7(490) <= '0';
partial_product_7(491) <= '0';
partial_product_7(492) <= '0';
partial_product_7(493) <= '0';
partial_product_7(494) <= '0';
partial_product_7(495) <= '0';
partial_product_7(496) <= '0';
partial_product_7(497) <= '0';
partial_product_7(498) <= '0';
partial_product_7(499) <= '0';
partial_product_7(500) <= '0';
partial_product_7(501) <= '0';
partial_product_7(502) <= '0';
partial_product_7(503) <= '0';
partial_product_7(504) <= '0';
partial_product_7(505) <= '0';
partial_product_7(506) <= '0';
partial_product_7(507) <= '0';
partial_product_7(508) <= '0';
partial_product_7(509) <= '0';
partial_product_7(510) <= '0';
partial_product_7(511) <= '0';
partial_product_7(512) <= '0';
partial_product_8(0) <= '0';
partial_product_8(1) <= '0';
partial_product_8(2) <= '0';
partial_product_8(3) <= '0';
partial_product_8(4) <= '0';
partial_product_8(5) <= '0';
partial_product_8(6) <= '0';
partial_product_8(7) <= '0';
partial_product_8(8) <= '0';
partial_product_8(9) <= '0';
partial_product_8(10) <= '0';
partial_product_8(11) <= '0';
partial_product_8(12) <= '0';
partial_product_8(13) <= '0';
partial_product_8(14) <= '0';
partial_product_8(15) <= '0';
partial_product_8(16) <= '0';
partial_product_8(17) <= '0';
partial_product_8(18) <= '0';
partial_product_8(19) <= '0';
partial_product_8(20) <= '0';
partial_product_8(21) <= '0';
partial_product_8(22) <= '0';
partial_product_8(23) <= '0';
partial_product_8(24) <= '0';
partial_product_8(25) <= '0';
partial_product_8(26) <= '0';
partial_product_8(27) <= '0';
partial_product_8(28) <= '0';
partial_product_8(29) <= '0';
partial_product_8(30) <= '0';
partial_product_8(31) <= '0';
partial_product_8(32) <= '0';
partial_product_8(33) <= '0';
partial_product_8(34) <= '0';
partial_product_8(35) <= '0';
partial_product_8(36) <= '0';
partial_product_8(37) <= '0';
partial_product_8(38) <= '0';
partial_product_8(39) <= '0';
partial_product_8(40) <= '0';
partial_product_8(41) <= '0';
partial_product_8(42) <= '0';
partial_product_8(43) <= '0';
partial_product_8(44) <= '0';
partial_product_8(45) <= '0';
partial_product_8(46) <= '0';
partial_product_8(47) <= '0';
partial_product_8(48) <= '0';
partial_product_8(49) <= '0';
partial_product_8(50) <= '0';
partial_product_8(51) <= '0';
partial_product_8(52) <= '0';
partial_product_8(53) <= '0';
partial_product_8(54) <= '0';
partial_product_8(55) <= '0';
partial_product_8(56) <= '0';
partial_product_8(57) <= '0';
partial_product_8(58) <= '0';
partial_product_8(59) <= '0';
partial_product_8(60) <= '0';
partial_product_8(61) <= '0';
partial_product_8(62) <= '0';
partial_product_8(63) <= '0';
partial_product_8(64) <= '0';
partial_product_8(65) <= '0';
partial_product_8(66) <= '0';
partial_product_8(67) <= '0';
partial_product_8(68) <= '0';
partial_product_8(69) <= '0';
partial_product_8(70) <= '0';
partial_product_8(71) <= '0';
partial_product_8(72) <= '0';
partial_product_8(73) <= '0';
partial_product_8(74) <= '0';
partial_product_8(75) <= '0';
partial_product_8(76) <= '0';
partial_product_8(77) <= '0';
partial_product_8(78) <= '0';
partial_product_8(79) <= '0';
partial_product_8(80) <= '0';
partial_product_8(81) <= '0';
partial_product_8(82) <= '0';
partial_product_8(83) <= '0';
partial_product_8(84) <= '0';
partial_product_8(85) <= temp_mult_25(85);
partial_product_8(86) <= temp_mult_25(86);
partial_product_8(87) <= temp_mult_25(87);
partial_product_8(88) <= temp_mult_25(88);
partial_product_8(89) <= temp_mult_25(89);
partial_product_8(90) <= temp_mult_25(90);
partial_product_8(91) <= temp_mult_25(91);
partial_product_8(92) <= temp_mult_25(92);
partial_product_8(93) <= temp_mult_25(93);
partial_product_8(94) <= temp_mult_25(94);
partial_product_8(95) <= temp_mult_25(95);
partial_product_8(96) <= temp_mult_25(96);
partial_product_8(97) <= temp_mult_25(97);
partial_product_8(98) <= temp_mult_25(98);
partial_product_8(99) <= temp_mult_25(99);
partial_product_8(100) <= temp_mult_25(100);
partial_product_8(101) <= temp_mult_25(101);
partial_product_8(102) <= temp_mult_25(102);
partial_product_8(103) <= temp_mult_25(103);
partial_product_8(104) <= temp_mult_25(104);
partial_product_8(105) <= temp_mult_25(105);
partial_product_8(106) <= temp_mult_25(106);
partial_product_8(107) <= temp_mult_25(107);
partial_product_8(108) <= temp_mult_25(108);
partial_product_8(109) <= temp_mult_25(109);
partial_product_8(110) <= temp_mult_25(110);
partial_product_8(111) <= temp_mult_25(111);
partial_product_8(112) <= temp_mult_25(112);
partial_product_8(113) <= temp_mult_25(113);
partial_product_8(114) <= temp_mult_25(114);
partial_product_8(115) <= temp_mult_25(115);
partial_product_8(116) <= temp_mult_25(116);
partial_product_8(117) <= temp_mult_25(117);
partial_product_8(118) <= temp_mult_25(118);
partial_product_8(119) <= temp_mult_25(119);
partial_product_8(120) <= temp_mult_25(120);
partial_product_8(121) <= temp_mult_25(121);
partial_product_8(122) <= temp_mult_25(122);
partial_product_8(123) <= temp_mult_25(123);
partial_product_8(124) <= temp_mult_25(124);
partial_product_8(125) <= temp_mult_25(125);
partial_product_8(126) <= temp_mult_31(126);
partial_product_8(127) <= temp_mult_31(127);
partial_product_8(128) <= temp_mult_31(128);
partial_product_8(129) <= temp_mult_31(129);
partial_product_8(130) <= temp_mult_31(130);
partial_product_8(131) <= temp_mult_31(131);
partial_product_8(132) <= temp_mult_31(132);
partial_product_8(133) <= temp_mult_31(133);
partial_product_8(134) <= temp_mult_31(134);
partial_product_8(135) <= temp_mult_31(135);
partial_product_8(136) <= temp_mult_31(136);
partial_product_8(137) <= temp_mult_31(137);
partial_product_8(138) <= temp_mult_31(138);
partial_product_8(139) <= temp_mult_31(139);
partial_product_8(140) <= temp_mult_31(140);
partial_product_8(141) <= temp_mult_31(141);
partial_product_8(142) <= temp_mult_31(142);
partial_product_8(143) <= temp_mult_31(143);
partial_product_8(144) <= temp_mult_31(144);
partial_product_8(145) <= temp_mult_31(145);
partial_product_8(146) <= temp_mult_31(146);
partial_product_8(147) <= temp_mult_31(147);
partial_product_8(148) <= temp_mult_31(148);
partial_product_8(149) <= temp_mult_31(149);
partial_product_8(150) <= temp_mult_31(150);
partial_product_8(151) <= temp_mult_31(151);
partial_product_8(152) <= temp_mult_31(152);
partial_product_8(153) <= temp_mult_31(153);
partial_product_8(154) <= temp_mult_31(154);
partial_product_8(155) <= temp_mult_31(155);
partial_product_8(156) <= temp_mult_31(156);
partial_product_8(157) <= temp_mult_31(157);
partial_product_8(158) <= temp_mult_31(158);
partial_product_8(159) <= temp_mult_31(159);
partial_product_8(160) <= temp_mult_31(160);
partial_product_8(161) <= temp_mult_31(161);
partial_product_8(162) <= temp_mult_31(162);
partial_product_8(163) <= temp_mult_31(163);
partial_product_8(164) <= temp_mult_31(164);
partial_product_8(165) <= temp_mult_31(165);
partial_product_8(166) <= temp_mult_31(166);
partial_product_8(167) <= temp_mult_37(167);
partial_product_8(168) <= temp_mult_37(168);
partial_product_8(169) <= temp_mult_37(169);
partial_product_8(170) <= temp_mult_37(170);
partial_product_8(171) <= temp_mult_37(171);
partial_product_8(172) <= temp_mult_37(172);
partial_product_8(173) <= temp_mult_37(173);
partial_product_8(174) <= temp_mult_37(174);
partial_product_8(175) <= temp_mult_37(175);
partial_product_8(176) <= temp_mult_37(176);
partial_product_8(177) <= temp_mult_37(177);
partial_product_8(178) <= temp_mult_37(178);
partial_product_8(179) <= temp_mult_37(179);
partial_product_8(180) <= temp_mult_37(180);
partial_product_8(181) <= temp_mult_37(181);
partial_product_8(182) <= temp_mult_37(182);
partial_product_8(183) <= temp_mult_37(183);
partial_product_8(184) <= temp_mult_37(184);
partial_product_8(185) <= temp_mult_37(185);
partial_product_8(186) <= temp_mult_37(186);
partial_product_8(187) <= temp_mult_37(187);
partial_product_8(188) <= temp_mult_37(188);
partial_product_8(189) <= temp_mult_37(189);
partial_product_8(190) <= temp_mult_37(190);
partial_product_8(191) <= temp_mult_37(191);
partial_product_8(192) <= temp_mult_37(192);
partial_product_8(193) <= temp_mult_37(193);
partial_product_8(194) <= temp_mult_37(194);
partial_product_8(195) <= temp_mult_37(195);
partial_product_8(196) <= temp_mult_37(196);
partial_product_8(197) <= temp_mult_37(197);
partial_product_8(198) <= temp_mult_37(198);
partial_product_8(199) <= temp_mult_37(199);
partial_product_8(200) <= temp_mult_37(200);
partial_product_8(201) <= temp_mult_37(201);
partial_product_8(202) <= temp_mult_37(202);
partial_product_8(203) <= temp_mult_37(203);
partial_product_8(204) <= temp_mult_37(204);
partial_product_8(205) <= temp_mult_37(205);
partial_product_8(206) <= temp_mult_37(206);
partial_product_8(207) <= temp_mult_37(207);
partial_product_8(208) <= temp_mult_104(208);
partial_product_8(209) <= temp_mult_104(209);
partial_product_8(210) <= temp_mult_104(210);
partial_product_8(211) <= temp_mult_104(211);
partial_product_8(212) <= temp_mult_104(212);
partial_product_8(213) <= temp_mult_104(213);
partial_product_8(214) <= temp_mult_104(214);
partial_product_8(215) <= temp_mult_104(215);
partial_product_8(216) <= temp_mult_104(216);
partial_product_8(217) <= temp_mult_104(217);
partial_product_8(218) <= temp_mult_104(218);
partial_product_8(219) <= temp_mult_104(219);
partial_product_8(220) <= temp_mult_104(220);
partial_product_8(221) <= temp_mult_104(221);
partial_product_8(222) <= temp_mult_104(222);
partial_product_8(223) <= temp_mult_104(223);
partial_product_8(224) <= temp_mult_104(224);
partial_product_8(225) <= temp_mult_104(225);
partial_product_8(226) <= temp_mult_104(226);
partial_product_8(227) <= temp_mult_104(227);
partial_product_8(228) <= temp_mult_104(228);
partial_product_8(229) <= temp_mult_104(229);
partial_product_8(230) <= temp_mult_104(230);
partial_product_8(231) <= temp_mult_104(231);
partial_product_8(232) <= temp_mult_104(232);
partial_product_8(233) <= temp_mult_104(233);
partial_product_8(234) <= temp_mult_104(234);
partial_product_8(235) <= temp_mult_104(235);
partial_product_8(236) <= temp_mult_104(236);
partial_product_8(237) <= temp_mult_104(237);
partial_product_8(238) <= temp_mult_104(238);
partial_product_8(239) <= temp_mult_104(239);
partial_product_8(240) <= temp_mult_104(240);
partial_product_8(241) <= temp_mult_104(241);
partial_product_8(242) <= temp_mult_104(242);
partial_product_8(243) <= temp_mult_104(243);
partial_product_8(244) <= temp_mult_104(244);
partial_product_8(245) <= temp_mult_104(245);
partial_product_8(246) <= temp_mult_104(246);
partial_product_8(247) <= temp_mult_104(247);
partial_product_8(248) <= temp_mult_104(248);
partial_product_8(249) <= temp_mult_113(249);
partial_product_8(250) <= temp_mult_113(250);
partial_product_8(251) <= temp_mult_113(251);
partial_product_8(252) <= temp_mult_113(252);
partial_product_8(253) <= temp_mult_113(253);
partial_product_8(254) <= temp_mult_113(254);
partial_product_8(255) <= temp_mult_113(255);
partial_product_8(256) <= temp_mult_113(256);
partial_product_8(257) <= temp_mult_113(257);
partial_product_8(258) <= temp_mult_113(258);
partial_product_8(259) <= temp_mult_113(259);
partial_product_8(260) <= temp_mult_113(260);
partial_product_8(261) <= temp_mult_113(261);
partial_product_8(262) <= temp_mult_113(262);
partial_product_8(263) <= temp_mult_113(263);
partial_product_8(264) <= temp_mult_113(264);
partial_product_8(265) <= temp_mult_113(265);
partial_product_8(266) <= temp_mult_113(266);
partial_product_8(267) <= temp_mult_113(267);
partial_product_8(268) <= temp_mult_113(268);
partial_product_8(269) <= temp_mult_113(269);
partial_product_8(270) <= temp_mult_113(270);
partial_product_8(271) <= temp_mult_113(271);
partial_product_8(272) <= temp_mult_113(272);
partial_product_8(273) <= temp_mult_113(273);
partial_product_8(274) <= temp_mult_113(274);
partial_product_8(275) <= temp_mult_113(275);
partial_product_8(276) <= temp_mult_113(276);
partial_product_8(277) <= temp_mult_113(277);
partial_product_8(278) <= temp_mult_113(278);
partial_product_8(279) <= temp_mult_113(279);
partial_product_8(280) <= temp_mult_113(280);
partial_product_8(281) <= temp_mult_113(281);
partial_product_8(282) <= temp_mult_113(282);
partial_product_8(283) <= temp_mult_113(283);
partial_product_8(284) <= temp_mult_113(284);
partial_product_8(285) <= temp_mult_113(285);
partial_product_8(286) <= temp_mult_113(286);
partial_product_8(287) <= temp_mult_113(287);
partial_product_8(288) <= temp_mult_113(288);
partial_product_8(289) <= temp_mult_113(289);
partial_product_8(290) <= temp_mult_130(290);
partial_product_8(291) <= temp_mult_130(291);
partial_product_8(292) <= temp_mult_130(292);
partial_product_8(293) <= temp_mult_130(293);
partial_product_8(294) <= temp_mult_130(294);
partial_product_8(295) <= temp_mult_130(295);
partial_product_8(296) <= temp_mult_130(296);
partial_product_8(297) <= temp_mult_130(297);
partial_product_8(298) <= temp_mult_130(298);
partial_product_8(299) <= temp_mult_130(299);
partial_product_8(300) <= temp_mult_130(300);
partial_product_8(301) <= temp_mult_130(301);
partial_product_8(302) <= temp_mult_130(302);
partial_product_8(303) <= temp_mult_130(303);
partial_product_8(304) <= temp_mult_130(304);
partial_product_8(305) <= temp_mult_130(305);
partial_product_8(306) <= temp_mult_130(306);
partial_product_8(307) <= temp_mult_130(307);
partial_product_8(308) <= temp_mult_130(308);
partial_product_8(309) <= temp_mult_130(309);
partial_product_8(310) <= temp_mult_130(310);
partial_product_8(311) <= temp_mult_130(311);
partial_product_8(312) <= temp_mult_130(312);
partial_product_8(313) <= temp_mult_130(313);
partial_product_8(314) <= temp_mult_130(314);
partial_product_8(315) <= temp_mult_130(315);
partial_product_8(316) <= temp_mult_130(316);
partial_product_8(317) <= temp_mult_130(317);
partial_product_8(318) <= temp_mult_130(318);
partial_product_8(319) <= temp_mult_130(319);
partial_product_8(320) <= temp_mult_130(320);
partial_product_8(321) <= temp_mult_130(321);
partial_product_8(322) <= temp_mult_130(322);
partial_product_8(323) <= temp_mult_130(323);
partial_product_8(324) <= temp_mult_130(324);
partial_product_8(325) <= temp_mult_130(325);
partial_product_8(326) <= temp_mult_130(326);
partial_product_8(327) <= temp_mult_130(327);
partial_product_8(328) <= temp_mult_130(328);
partial_product_8(329) <= temp_mult_130(329);
partial_product_8(330) <= temp_mult_130(330);
partial_product_8(331) <= temp_mult_136(331);
partial_product_8(332) <= temp_mult_136(332);
partial_product_8(333) <= temp_mult_136(333);
partial_product_8(334) <= temp_mult_136(334);
partial_product_8(335) <= temp_mult_136(335);
partial_product_8(336) <= temp_mult_136(336);
partial_product_8(337) <= temp_mult_136(337);
partial_product_8(338) <= temp_mult_136(338);
partial_product_8(339) <= temp_mult_136(339);
partial_product_8(340) <= temp_mult_136(340);
partial_product_8(341) <= temp_mult_136(341);
partial_product_8(342) <= temp_mult_136(342);
partial_product_8(343) <= temp_mult_136(343);
partial_product_8(344) <= temp_mult_136(344);
partial_product_8(345) <= temp_mult_136(345);
partial_product_8(346) <= temp_mult_136(346);
partial_product_8(347) <= temp_mult_136(347);
partial_product_8(348) <= temp_mult_136(348);
partial_product_8(349) <= temp_mult_136(349);
partial_product_8(350) <= temp_mult_136(350);
partial_product_8(351) <= temp_mult_136(351);
partial_product_8(352) <= temp_mult_136(352);
partial_product_8(353) <= temp_mult_136(353);
partial_product_8(354) <= temp_mult_136(354);
partial_product_8(355) <= temp_mult_136(355);
partial_product_8(356) <= temp_mult_136(356);
partial_product_8(357) <= temp_mult_136(357);
partial_product_8(358) <= temp_mult_136(358);
partial_product_8(359) <= temp_mult_136(359);
partial_product_8(360) <= temp_mult_136(360);
partial_product_8(361) <= temp_mult_136(361);
partial_product_8(362) <= temp_mult_136(362);
partial_product_8(363) <= temp_mult_136(363);
partial_product_8(364) <= temp_mult_136(364);
partial_product_8(365) <= temp_mult_136(365);
partial_product_8(366) <= temp_mult_136(366);
partial_product_8(367) <= temp_mult_136(367);
partial_product_8(368) <= temp_mult_136(368);
partial_product_8(369) <= temp_mult_136(369);
partial_product_8(370) <= temp_mult_136(370);
partial_product_8(371) <= temp_mult_136(371);
partial_product_8(372) <= temp_mult_142(372);
partial_product_8(373) <= temp_mult_142(373);
partial_product_8(374) <= temp_mult_142(374);
partial_product_8(375) <= temp_mult_142(375);
partial_product_8(376) <= temp_mult_142(376);
partial_product_8(377) <= temp_mult_142(377);
partial_product_8(378) <= temp_mult_142(378);
partial_product_8(379) <= temp_mult_142(379);
partial_product_8(380) <= temp_mult_142(380);
partial_product_8(381) <= temp_mult_142(381);
partial_product_8(382) <= temp_mult_142(382);
partial_product_8(383) <= temp_mult_142(383);
partial_product_8(384) <= temp_mult_142(384);
partial_product_8(385) <= temp_mult_142(385);
partial_product_8(386) <= temp_mult_142(386);
partial_product_8(387) <= temp_mult_142(387);
partial_product_8(388) <= temp_mult_142(388);
partial_product_8(389) <= temp_mult_142(389);
partial_product_8(390) <= temp_mult_142(390);
partial_product_8(391) <= temp_mult_142(391);
partial_product_8(392) <= temp_mult_142(392);
partial_product_8(393) <= temp_mult_142(393);
partial_product_8(394) <= temp_mult_142(394);
partial_product_8(395) <= temp_mult_142(395);
partial_product_8(396) <= temp_mult_142(396);
partial_product_8(397) <= temp_mult_142(397);
partial_product_8(398) <= temp_mult_142(398);
partial_product_8(399) <= temp_mult_142(399);
partial_product_8(400) <= temp_mult_142(400);
partial_product_8(401) <= temp_mult_142(401);
partial_product_8(402) <= temp_mult_142(402);
partial_product_8(403) <= temp_mult_142(403);
partial_product_8(404) <= temp_mult_142(404);
partial_product_8(405) <= temp_mult_142(405);
partial_product_8(406) <= temp_mult_142(406);
partial_product_8(407) <= temp_mult_142(407);
partial_product_8(408) <= temp_mult_142(408);
partial_product_8(409) <= temp_mult_142(409);
partial_product_8(410) <= temp_mult_142(410);
partial_product_8(411) <= temp_mult_142(411);
partial_product_8(412) <= temp_mult_142(412);
partial_product_8(413) <= '0';
partial_product_8(414) <= '0';
partial_product_8(415) <= '0';
partial_product_8(416) <= '0';
partial_product_8(417) <= '0';
partial_product_8(418) <= '0';
partial_product_8(419) <= '0';
partial_product_8(420) <= '0';
partial_product_8(421) <= '0';
partial_product_8(422) <= '0';
partial_product_8(423) <= '0';
partial_product_8(424) <= '0';
partial_product_8(425) <= '0';
partial_product_8(426) <= '0';
partial_product_8(427) <= '0';
partial_product_8(428) <= '0';
partial_product_8(429) <= '0';
partial_product_8(430) <= '0';
partial_product_8(431) <= '0';
partial_product_8(432) <= '0';
partial_product_8(433) <= '0';
partial_product_8(434) <= '0';
partial_product_8(435) <= '0';
partial_product_8(436) <= '0';
partial_product_8(437) <= '0';
partial_product_8(438) <= '0';
partial_product_8(439) <= '0';
partial_product_8(440) <= '0';
partial_product_8(441) <= '0';
partial_product_8(442) <= '0';
partial_product_8(443) <= '0';
partial_product_8(444) <= '0';
partial_product_8(445) <= '0';
partial_product_8(446) <= '0';
partial_product_8(447) <= '0';
partial_product_8(448) <= '0';
partial_product_8(449) <= '0';
partial_product_8(450) <= '0';
partial_product_8(451) <= '0';
partial_product_8(452) <= '0';
partial_product_8(453) <= '0';
partial_product_8(454) <= '0';
partial_product_8(455) <= '0';
partial_product_8(456) <= '0';
partial_product_8(457) <= '0';
partial_product_8(458) <= '0';
partial_product_8(459) <= '0';
partial_product_8(460) <= '0';
partial_product_8(461) <= '0';
partial_product_8(462) <= '0';
partial_product_8(463) <= '0';
partial_product_8(464) <= '0';
partial_product_8(465) <= '0';
partial_product_8(466) <= '0';
partial_product_8(467) <= '0';
partial_product_8(468) <= '0';
partial_product_8(469) <= '0';
partial_product_8(470) <= '0';
partial_product_8(471) <= '0';
partial_product_8(472) <= '0';
partial_product_8(473) <= '0';
partial_product_8(474) <= '0';
partial_product_8(475) <= '0';
partial_product_8(476) <= '0';
partial_product_8(477) <= '0';
partial_product_8(478) <= '0';
partial_product_8(479) <= '0';
partial_product_8(480) <= '0';
partial_product_8(481) <= '0';
partial_product_8(482) <= '0';
partial_product_8(483) <= '0';
partial_product_8(484) <= '0';
partial_product_8(485) <= '0';
partial_product_8(486) <= '0';
partial_product_8(487) <= '0';
partial_product_8(488) <= '0';
partial_product_8(489) <= '0';
partial_product_8(490) <= '0';
partial_product_8(491) <= '0';
partial_product_8(492) <= '0';
partial_product_8(493) <= '0';
partial_product_8(494) <= '0';
partial_product_8(495) <= '0';
partial_product_8(496) <= '0';
partial_product_8(497) <= '0';
partial_product_8(498) <= '0';
partial_product_8(499) <= '0';
partial_product_8(500) <= '0';
partial_product_8(501) <= '0';
partial_product_8(502) <= '0';
partial_product_8(503) <= '0';
partial_product_8(504) <= '0';
partial_product_8(505) <= '0';
partial_product_8(506) <= '0';
partial_product_8(507) <= '0';
partial_product_8(508) <= '0';
partial_product_8(509) <= '0';
partial_product_8(510) <= '0';
partial_product_8(511) <= '0';
partial_product_8(512) <= '0';
partial_product_9(0) <= '0';
partial_product_9(1) <= '0';
partial_product_9(2) <= '0';
partial_product_9(3) <= '0';
partial_product_9(4) <= '0';
partial_product_9(5) <= '0';
partial_product_9(6) <= '0';
partial_product_9(7) <= '0';
partial_product_9(8) <= '0';
partial_product_9(9) <= '0';
partial_product_9(10) <= '0';
partial_product_9(11) <= '0';
partial_product_9(12) <= '0';
partial_product_9(13) <= '0';
partial_product_9(14) <= '0';
partial_product_9(15) <= '0';
partial_product_9(16) <= '0';
partial_product_9(17) <= '0';
partial_product_9(18) <= '0';
partial_product_9(19) <= '0';
partial_product_9(20) <= '0';
partial_product_9(21) <= '0';
partial_product_9(22) <= '0';
partial_product_9(23) <= '0';
partial_product_9(24) <= '0';
partial_product_9(25) <= '0';
partial_product_9(26) <= '0';
partial_product_9(27) <= '0';
partial_product_9(28) <= '0';
partial_product_9(29) <= '0';
partial_product_9(30) <= '0';
partial_product_9(31) <= '0';
partial_product_9(32) <= '0';
partial_product_9(33) <= '0';
partial_product_9(34) <= '0';
partial_product_9(35) <= '0';
partial_product_9(36) <= '0';
partial_product_9(37) <= '0';
partial_product_9(38) <= '0';
partial_product_9(39) <= '0';
partial_product_9(40) <= '0';
partial_product_9(41) <= '0';
partial_product_9(42) <= '0';
partial_product_9(43) <= '0';
partial_product_9(44) <= '0';
partial_product_9(45) <= '0';
partial_product_9(46) <= '0';
partial_product_9(47) <= '0';
partial_product_9(48) <= '0';
partial_product_9(49) <= '0';
partial_product_9(50) <= '0';
partial_product_9(51) <= '0';
partial_product_9(52) <= '0';
partial_product_9(53) <= '0';
partial_product_9(54) <= '0';
partial_product_9(55) <= '0';
partial_product_9(56) <= '0';
partial_product_9(57) <= '0';
partial_product_9(58) <= '0';
partial_product_9(59) <= '0';
partial_product_9(60) <= '0';
partial_product_9(61) <= '0';
partial_product_9(62) <= '0';
partial_product_9(63) <= '0';
partial_product_9(64) <= '0';
partial_product_9(65) <= '0';
partial_product_9(66) <= '0';
partial_product_9(67) <= '0';
partial_product_9(68) <= '0';
partial_product_9(69) <= '0';
partial_product_9(70) <= '0';
partial_product_9(71) <= '0';
partial_product_9(72) <= '0';
partial_product_9(73) <= '0';
partial_product_9(74) <= '0';
partial_product_9(75) <= '0';
partial_product_9(76) <= '0';
partial_product_9(77) <= '0';
partial_product_9(78) <= '0';
partial_product_9(79) <= '0';
partial_product_9(80) <= '0';
partial_product_9(81) <= '0';
partial_product_9(82) <= '0';
partial_product_9(83) <= '0';
partial_product_9(84) <= '0';
partial_product_9(85) <= '0';
partial_product_9(86) <= '0';
partial_product_9(87) <= '0';
partial_product_9(88) <= '0';
partial_product_9(89) <= '0';
partial_product_9(90) <= '0';
partial_product_9(91) <= '0';
partial_product_9(92) <= '0';
partial_product_9(93) <= '0';
partial_product_9(94) <= '0';
partial_product_9(95) <= '0';
partial_product_9(96) <= temp_mult_4(96);
partial_product_9(97) <= temp_mult_4(97);
partial_product_9(98) <= temp_mult_4(98);
partial_product_9(99) <= temp_mult_4(99);
partial_product_9(100) <= temp_mult_4(100);
partial_product_9(101) <= temp_mult_4(101);
partial_product_9(102) <= temp_mult_4(102);
partial_product_9(103) <= temp_mult_4(103);
partial_product_9(104) <= temp_mult_4(104);
partial_product_9(105) <= temp_mult_4(105);
partial_product_9(106) <= temp_mult_4(106);
partial_product_9(107) <= temp_mult_4(107);
partial_product_9(108) <= temp_mult_4(108);
partial_product_9(109) <= temp_mult_4(109);
partial_product_9(110) <= temp_mult_4(110);
partial_product_9(111) <= temp_mult_4(111);
partial_product_9(112) <= temp_mult_4(112);
partial_product_9(113) <= temp_mult_4(113);
partial_product_9(114) <= temp_mult_4(114);
partial_product_9(115) <= temp_mult_4(115);
partial_product_9(116) <= temp_mult_4(116);
partial_product_9(117) <= temp_mult_4(117);
partial_product_9(118) <= temp_mult_4(118);
partial_product_9(119) <= temp_mult_4(119);
partial_product_9(120) <= temp_mult_4(120);
partial_product_9(121) <= temp_mult_4(121);
partial_product_9(122) <= temp_mult_4(122);
partial_product_9(123) <= temp_mult_4(123);
partial_product_9(124) <= temp_mult_4(124);
partial_product_9(125) <= temp_mult_4(125);
partial_product_9(126) <= temp_mult_4(126);
partial_product_9(127) <= temp_mult_4(127);
partial_product_9(128) <= temp_mult_4(128);
partial_product_9(129) <= temp_mult_4(129);
partial_product_9(130) <= temp_mult_4(130);
partial_product_9(131) <= temp_mult_4(131);
partial_product_9(132) <= temp_mult_4(132);
partial_product_9(133) <= temp_mult_4(133);
partial_product_9(134) <= temp_mult_4(134);
partial_product_9(135) <= temp_mult_4(135);
partial_product_9(136) <= temp_mult_4(136);
partial_product_9(137) <= temp_mult_41(137);
partial_product_9(138) <= temp_mult_41(138);
partial_product_9(139) <= temp_mult_41(139);
partial_product_9(140) <= temp_mult_41(140);
partial_product_9(141) <= temp_mult_41(141);
partial_product_9(142) <= temp_mult_41(142);
partial_product_9(143) <= temp_mult_41(143);
partial_product_9(144) <= temp_mult_41(144);
partial_product_9(145) <= temp_mult_41(145);
partial_product_9(146) <= temp_mult_41(146);
partial_product_9(147) <= temp_mult_41(147);
partial_product_9(148) <= temp_mult_41(148);
partial_product_9(149) <= temp_mult_41(149);
partial_product_9(150) <= temp_mult_41(150);
partial_product_9(151) <= temp_mult_41(151);
partial_product_9(152) <= temp_mult_41(152);
partial_product_9(153) <= temp_mult_41(153);
partial_product_9(154) <= temp_mult_41(154);
partial_product_9(155) <= temp_mult_41(155);
partial_product_9(156) <= temp_mult_41(156);
partial_product_9(157) <= temp_mult_41(157);
partial_product_9(158) <= temp_mult_41(158);
partial_product_9(159) <= temp_mult_41(159);
partial_product_9(160) <= temp_mult_41(160);
partial_product_9(161) <= temp_mult_41(161);
partial_product_9(162) <= temp_mult_41(162);
partial_product_9(163) <= temp_mult_41(163);
partial_product_9(164) <= temp_mult_41(164);
partial_product_9(165) <= temp_mult_41(165);
partial_product_9(166) <= temp_mult_41(166);
partial_product_9(167) <= temp_mult_41(167);
partial_product_9(168) <= temp_mult_41(168);
partial_product_9(169) <= temp_mult_41(169);
partial_product_9(170) <= temp_mult_41(170);
partial_product_9(171) <= temp_mult_41(171);
partial_product_9(172) <= temp_mult_41(172);
partial_product_9(173) <= temp_mult_41(173);
partial_product_9(174) <= temp_mult_41(174);
partial_product_9(175) <= temp_mult_41(175);
partial_product_9(176) <= temp_mult_41(176);
partial_product_9(177) <= temp_mult_41(177);
partial_product_9(178) <= temp_mult_50(178);
partial_product_9(179) <= temp_mult_50(179);
partial_product_9(180) <= temp_mult_50(180);
partial_product_9(181) <= temp_mult_50(181);
partial_product_9(182) <= temp_mult_50(182);
partial_product_9(183) <= temp_mult_50(183);
partial_product_9(184) <= temp_mult_50(184);
partial_product_9(185) <= temp_mult_50(185);
partial_product_9(186) <= temp_mult_50(186);
partial_product_9(187) <= temp_mult_50(187);
partial_product_9(188) <= temp_mult_50(188);
partial_product_9(189) <= temp_mult_50(189);
partial_product_9(190) <= temp_mult_50(190);
partial_product_9(191) <= temp_mult_50(191);
partial_product_9(192) <= temp_mult_50(192);
partial_product_9(193) <= temp_mult_50(193);
partial_product_9(194) <= temp_mult_50(194);
partial_product_9(195) <= temp_mult_50(195);
partial_product_9(196) <= temp_mult_50(196);
partial_product_9(197) <= temp_mult_50(197);
partial_product_9(198) <= temp_mult_50(198);
partial_product_9(199) <= temp_mult_50(199);
partial_product_9(200) <= temp_mult_50(200);
partial_product_9(201) <= temp_mult_50(201);
partial_product_9(202) <= temp_mult_50(202);
partial_product_9(203) <= temp_mult_50(203);
partial_product_9(204) <= temp_mult_50(204);
partial_product_9(205) <= temp_mult_50(205);
partial_product_9(206) <= temp_mult_50(206);
partial_product_9(207) <= temp_mult_50(207);
partial_product_9(208) <= temp_mult_50(208);
partial_product_9(209) <= temp_mult_50(209);
partial_product_9(210) <= temp_mult_50(210);
partial_product_9(211) <= temp_mult_50(211);
partial_product_9(212) <= temp_mult_50(212);
partial_product_9(213) <= temp_mult_50(213);
partial_product_9(214) <= temp_mult_50(214);
partial_product_9(215) <= temp_mult_50(215);
partial_product_9(216) <= temp_mult_50(216);
partial_product_9(217) <= temp_mult_50(217);
partial_product_9(218) <= temp_mult_50(218);
partial_product_9(219) <= temp_mult_59(219);
partial_product_9(220) <= temp_mult_59(220);
partial_product_9(221) <= temp_mult_59(221);
partial_product_9(222) <= temp_mult_59(222);
partial_product_9(223) <= temp_mult_59(223);
partial_product_9(224) <= temp_mult_59(224);
partial_product_9(225) <= temp_mult_59(225);
partial_product_9(226) <= temp_mult_59(226);
partial_product_9(227) <= temp_mult_59(227);
partial_product_9(228) <= temp_mult_59(228);
partial_product_9(229) <= temp_mult_59(229);
partial_product_9(230) <= temp_mult_59(230);
partial_product_9(231) <= temp_mult_59(231);
partial_product_9(232) <= temp_mult_59(232);
partial_product_9(233) <= temp_mult_59(233);
partial_product_9(234) <= temp_mult_59(234);
partial_product_9(235) <= temp_mult_59(235);
partial_product_9(236) <= temp_mult_59(236);
partial_product_9(237) <= temp_mult_59(237);
partial_product_9(238) <= temp_mult_59(238);
partial_product_9(239) <= temp_mult_59(239);
partial_product_9(240) <= temp_mult_59(240);
partial_product_9(241) <= temp_mult_59(241);
partial_product_9(242) <= temp_mult_59(242);
partial_product_9(243) <= temp_mult_59(243);
partial_product_9(244) <= temp_mult_59(244);
partial_product_9(245) <= temp_mult_59(245);
partial_product_9(246) <= temp_mult_59(246);
partial_product_9(247) <= temp_mult_59(247);
partial_product_9(248) <= temp_mult_59(248);
partial_product_9(249) <= temp_mult_59(249);
partial_product_9(250) <= temp_mult_59(250);
partial_product_9(251) <= temp_mult_59(251);
partial_product_9(252) <= temp_mult_59(252);
partial_product_9(253) <= temp_mult_59(253);
partial_product_9(254) <= temp_mult_59(254);
partial_product_9(255) <= temp_mult_59(255);
partial_product_9(256) <= temp_mult_59(256);
partial_product_9(257) <= temp_mult_59(257);
partial_product_9(258) <= temp_mult_59(258);
partial_product_9(259) <= temp_mult_59(259);
partial_product_9(260) <= temp_mult_68(260);
partial_product_9(261) <= temp_mult_68(261);
partial_product_9(262) <= temp_mult_68(262);
partial_product_9(263) <= temp_mult_68(263);
partial_product_9(264) <= temp_mult_68(264);
partial_product_9(265) <= temp_mult_68(265);
partial_product_9(266) <= temp_mult_68(266);
partial_product_9(267) <= temp_mult_68(267);
partial_product_9(268) <= temp_mult_68(268);
partial_product_9(269) <= temp_mult_68(269);
partial_product_9(270) <= temp_mult_68(270);
partial_product_9(271) <= temp_mult_68(271);
partial_product_9(272) <= temp_mult_68(272);
partial_product_9(273) <= temp_mult_68(273);
partial_product_9(274) <= temp_mult_68(274);
partial_product_9(275) <= temp_mult_68(275);
partial_product_9(276) <= temp_mult_68(276);
partial_product_9(277) <= temp_mult_68(277);
partial_product_9(278) <= temp_mult_68(278);
partial_product_9(279) <= temp_mult_68(279);
partial_product_9(280) <= temp_mult_68(280);
partial_product_9(281) <= temp_mult_68(281);
partial_product_9(282) <= temp_mult_68(282);
partial_product_9(283) <= temp_mult_68(283);
partial_product_9(284) <= temp_mult_68(284);
partial_product_9(285) <= temp_mult_68(285);
partial_product_9(286) <= temp_mult_68(286);
partial_product_9(287) <= temp_mult_68(287);
partial_product_9(288) <= temp_mult_68(288);
partial_product_9(289) <= temp_mult_68(289);
partial_product_9(290) <= temp_mult_68(290);
partial_product_9(291) <= temp_mult_68(291);
partial_product_9(292) <= temp_mult_68(292);
partial_product_9(293) <= temp_mult_68(293);
partial_product_9(294) <= temp_mult_68(294);
partial_product_9(295) <= temp_mult_68(295);
partial_product_9(296) <= temp_mult_68(296);
partial_product_9(297) <= temp_mult_68(297);
partial_product_9(298) <= temp_mult_68(298);
partial_product_9(299) <= temp_mult_68(299);
partial_product_9(300) <= temp_mult_68(300);
partial_product_9(301) <= temp_mult_77(301);
partial_product_9(302) <= temp_mult_77(302);
partial_product_9(303) <= temp_mult_77(303);
partial_product_9(304) <= temp_mult_77(304);
partial_product_9(305) <= temp_mult_77(305);
partial_product_9(306) <= temp_mult_77(306);
partial_product_9(307) <= temp_mult_77(307);
partial_product_9(308) <= temp_mult_77(308);
partial_product_9(309) <= temp_mult_77(309);
partial_product_9(310) <= temp_mult_77(310);
partial_product_9(311) <= temp_mult_77(311);
partial_product_9(312) <= temp_mult_77(312);
partial_product_9(313) <= temp_mult_77(313);
partial_product_9(314) <= temp_mult_77(314);
partial_product_9(315) <= temp_mult_77(315);
partial_product_9(316) <= temp_mult_77(316);
partial_product_9(317) <= temp_mult_77(317);
partial_product_9(318) <= temp_mult_77(318);
partial_product_9(319) <= temp_mult_77(319);
partial_product_9(320) <= temp_mult_77(320);
partial_product_9(321) <= temp_mult_77(321);
partial_product_9(322) <= temp_mult_77(322);
partial_product_9(323) <= temp_mult_77(323);
partial_product_9(324) <= temp_mult_77(324);
partial_product_9(325) <= temp_mult_77(325);
partial_product_9(326) <= temp_mult_77(326);
partial_product_9(327) <= temp_mult_77(327);
partial_product_9(328) <= temp_mult_77(328);
partial_product_9(329) <= temp_mult_77(329);
partial_product_9(330) <= temp_mult_77(330);
partial_product_9(331) <= temp_mult_77(331);
partial_product_9(332) <= temp_mult_77(332);
partial_product_9(333) <= temp_mult_77(333);
partial_product_9(334) <= temp_mult_77(334);
partial_product_9(335) <= temp_mult_77(335);
partial_product_9(336) <= temp_mult_77(336);
partial_product_9(337) <= temp_mult_77(337);
partial_product_9(338) <= temp_mult_77(338);
partial_product_9(339) <= temp_mult_77(339);
partial_product_9(340) <= temp_mult_77(340);
partial_product_9(341) <= temp_mult_77(341);
partial_product_9(342) <= '0';
partial_product_9(343) <= '0';
partial_product_9(344) <= '0';
partial_product_9(345) <= '0';
partial_product_9(346) <= '0';
partial_product_9(347) <= '0';
partial_product_9(348) <= temp_mult_141(348);
partial_product_9(349) <= temp_mult_141(349);
partial_product_9(350) <= temp_mult_141(350);
partial_product_9(351) <= temp_mult_141(351);
partial_product_9(352) <= temp_mult_141(352);
partial_product_9(353) <= temp_mult_141(353);
partial_product_9(354) <= temp_mult_141(354);
partial_product_9(355) <= temp_mult_141(355);
partial_product_9(356) <= temp_mult_141(356);
partial_product_9(357) <= temp_mult_141(357);
partial_product_9(358) <= temp_mult_141(358);
partial_product_9(359) <= temp_mult_141(359);
partial_product_9(360) <= temp_mult_141(360);
partial_product_9(361) <= temp_mult_141(361);
partial_product_9(362) <= temp_mult_141(362);
partial_product_9(363) <= temp_mult_141(363);
partial_product_9(364) <= temp_mult_141(364);
partial_product_9(365) <= temp_mult_141(365);
partial_product_9(366) <= temp_mult_141(366);
partial_product_9(367) <= temp_mult_141(367);
partial_product_9(368) <= temp_mult_141(368);
partial_product_9(369) <= temp_mult_141(369);
partial_product_9(370) <= temp_mult_141(370);
partial_product_9(371) <= temp_mult_141(371);
partial_product_9(372) <= temp_mult_141(372);
partial_product_9(373) <= temp_mult_141(373);
partial_product_9(374) <= temp_mult_141(374);
partial_product_9(375) <= temp_mult_141(375);
partial_product_9(376) <= temp_mult_141(376);
partial_product_9(377) <= temp_mult_141(377);
partial_product_9(378) <= temp_mult_141(378);
partial_product_9(379) <= temp_mult_141(379);
partial_product_9(380) <= temp_mult_141(380);
partial_product_9(381) <= temp_mult_141(381);
partial_product_9(382) <= temp_mult_141(382);
partial_product_9(383) <= temp_mult_141(383);
partial_product_9(384) <= temp_mult_141(384);
partial_product_9(385) <= temp_mult_141(385);
partial_product_9(386) <= temp_mult_141(386);
partial_product_9(387) <= temp_mult_141(387);
partial_product_9(388) <= temp_mult_141(388);
partial_product_9(389) <= temp_mult_147(389);
partial_product_9(390) <= temp_mult_147(390);
partial_product_9(391) <= temp_mult_147(391);
partial_product_9(392) <= temp_mult_147(392);
partial_product_9(393) <= temp_mult_147(393);
partial_product_9(394) <= temp_mult_147(394);
partial_product_9(395) <= temp_mult_147(395);
partial_product_9(396) <= temp_mult_147(396);
partial_product_9(397) <= temp_mult_147(397);
partial_product_9(398) <= temp_mult_147(398);
partial_product_9(399) <= temp_mult_147(399);
partial_product_9(400) <= temp_mult_147(400);
partial_product_9(401) <= temp_mult_147(401);
partial_product_9(402) <= temp_mult_147(402);
partial_product_9(403) <= temp_mult_147(403);
partial_product_9(404) <= temp_mult_147(404);
partial_product_9(405) <= temp_mult_147(405);
partial_product_9(406) <= temp_mult_147(406);
partial_product_9(407) <= temp_mult_147(407);
partial_product_9(408) <= temp_mult_147(408);
partial_product_9(409) <= temp_mult_147(409);
partial_product_9(410) <= temp_mult_147(410);
partial_product_9(411) <= temp_mult_147(411);
partial_product_9(412) <= temp_mult_147(412);
partial_product_9(413) <= temp_mult_147(413);
partial_product_9(414) <= temp_mult_147(414);
partial_product_9(415) <= temp_mult_147(415);
partial_product_9(416) <= temp_mult_147(416);
partial_product_9(417) <= temp_mult_147(417);
partial_product_9(418) <= temp_mult_147(418);
partial_product_9(419) <= temp_mult_147(419);
partial_product_9(420) <= temp_mult_147(420);
partial_product_9(421) <= temp_mult_147(421);
partial_product_9(422) <= temp_mult_147(422);
partial_product_9(423) <= temp_mult_147(423);
partial_product_9(424) <= temp_mult_147(424);
partial_product_9(425) <= temp_mult_147(425);
partial_product_9(426) <= temp_mult_147(426);
partial_product_9(427) <= temp_mult_147(427);
partial_product_9(428) <= temp_mult_147(428);
partial_product_9(429) <= temp_mult_147(429);
partial_product_9(430) <= '0';
partial_product_9(431) <= '0';
partial_product_9(432) <= '0';
partial_product_9(433) <= '0';
partial_product_9(434) <= '0';
partial_product_9(435) <= '0';
partial_product_9(436) <= '0';
partial_product_9(437) <= '0';
partial_product_9(438) <= '0';
partial_product_9(439) <= '0';
partial_product_9(440) <= '0';
partial_product_9(441) <= '0';
partial_product_9(442) <= '0';
partial_product_9(443) <= '0';
partial_product_9(444) <= '0';
partial_product_9(445) <= '0';
partial_product_9(446) <= '0';
partial_product_9(447) <= '0';
partial_product_9(448) <= '0';
partial_product_9(449) <= '0';
partial_product_9(450) <= '0';
partial_product_9(451) <= '0';
partial_product_9(452) <= '0';
partial_product_9(453) <= '0';
partial_product_9(454) <= '0';
partial_product_9(455) <= '0';
partial_product_9(456) <= '0';
partial_product_9(457) <= '0';
partial_product_9(458) <= '0';
partial_product_9(459) <= '0';
partial_product_9(460) <= '0';
partial_product_9(461) <= '0';
partial_product_9(462) <= '0';
partial_product_9(463) <= '0';
partial_product_9(464) <= '0';
partial_product_9(465) <= '0';
partial_product_9(466) <= '0';
partial_product_9(467) <= '0';
partial_product_9(468) <= '0';
partial_product_9(469) <= '0';
partial_product_9(470) <= '0';
partial_product_9(471) <= '0';
partial_product_9(472) <= '0';
partial_product_9(473) <= '0';
partial_product_9(474) <= '0';
partial_product_9(475) <= '0';
partial_product_9(476) <= '0';
partial_product_9(477) <= '0';
partial_product_9(478) <= '0';
partial_product_9(479) <= '0';
partial_product_9(480) <= '0';
partial_product_9(481) <= '0';
partial_product_9(482) <= '0';
partial_product_9(483) <= '0';
partial_product_9(484) <= '0';
partial_product_9(485) <= '0';
partial_product_9(486) <= '0';
partial_product_9(487) <= '0';
partial_product_9(488) <= '0';
partial_product_9(489) <= '0';
partial_product_9(490) <= '0';
partial_product_9(491) <= '0';
partial_product_9(492) <= '0';
partial_product_9(493) <= '0';
partial_product_9(494) <= '0';
partial_product_9(495) <= '0';
partial_product_9(496) <= '0';
partial_product_9(497) <= '0';
partial_product_9(498) <= '0';
partial_product_9(499) <= '0';
partial_product_9(500) <= '0';
partial_product_9(501) <= '0';
partial_product_9(502) <= '0';
partial_product_9(503) <= '0';
partial_product_9(504) <= '0';
partial_product_9(505) <= '0';
partial_product_9(506) <= '0';
partial_product_9(507) <= '0';
partial_product_9(508) <= '0';
partial_product_9(509) <= '0';
partial_product_9(510) <= '0';
partial_product_9(511) <= '0';
partial_product_9(512) <= '0';
partial_product_10(0) <= '0';
partial_product_10(1) <= '0';
partial_product_10(2) <= '0';
partial_product_10(3) <= '0';
partial_product_10(4) <= '0';
partial_product_10(5) <= '0';
partial_product_10(6) <= '0';
partial_product_10(7) <= '0';
partial_product_10(8) <= '0';
partial_product_10(9) <= '0';
partial_product_10(10) <= '0';
partial_product_10(11) <= '0';
partial_product_10(12) <= '0';
partial_product_10(13) <= '0';
partial_product_10(14) <= '0';
partial_product_10(15) <= '0';
partial_product_10(16) <= '0';
partial_product_10(17) <= '0';
partial_product_10(18) <= '0';
partial_product_10(19) <= '0';
partial_product_10(20) <= '0';
partial_product_10(21) <= '0';
partial_product_10(22) <= '0';
partial_product_10(23) <= '0';
partial_product_10(24) <= '0';
partial_product_10(25) <= '0';
partial_product_10(26) <= '0';
partial_product_10(27) <= '0';
partial_product_10(28) <= '0';
partial_product_10(29) <= '0';
partial_product_10(30) <= '0';
partial_product_10(31) <= '0';
partial_product_10(32) <= '0';
partial_product_10(33) <= '0';
partial_product_10(34) <= '0';
partial_product_10(35) <= '0';
partial_product_10(36) <= '0';
partial_product_10(37) <= '0';
partial_product_10(38) <= '0';
partial_product_10(39) <= '0';
partial_product_10(40) <= '0';
partial_product_10(41) <= '0';
partial_product_10(42) <= '0';
partial_product_10(43) <= '0';
partial_product_10(44) <= '0';
partial_product_10(45) <= '0';
partial_product_10(46) <= '0';
partial_product_10(47) <= '0';
partial_product_10(48) <= '0';
partial_product_10(49) <= '0';
partial_product_10(50) <= '0';
partial_product_10(51) <= '0';
partial_product_10(52) <= '0';
partial_product_10(53) <= '0';
partial_product_10(54) <= '0';
partial_product_10(55) <= '0';
partial_product_10(56) <= '0';
partial_product_10(57) <= '0';
partial_product_10(58) <= '0';
partial_product_10(59) <= '0';
partial_product_10(60) <= '0';
partial_product_10(61) <= '0';
partial_product_10(62) <= '0';
partial_product_10(63) <= '0';
partial_product_10(64) <= '0';
partial_product_10(65) <= '0';
partial_product_10(66) <= '0';
partial_product_10(67) <= '0';
partial_product_10(68) <= '0';
partial_product_10(69) <= '0';
partial_product_10(70) <= '0';
partial_product_10(71) <= '0';
partial_product_10(72) <= '0';
partial_product_10(73) <= '0';
partial_product_10(74) <= '0';
partial_product_10(75) <= '0';
partial_product_10(76) <= '0';
partial_product_10(77) <= '0';
partial_product_10(78) <= '0';
partial_product_10(79) <= '0';
partial_product_10(80) <= '0';
partial_product_10(81) <= '0';
partial_product_10(82) <= '0';
partial_product_10(83) <= '0';
partial_product_10(84) <= '0';
partial_product_10(85) <= '0';
partial_product_10(86) <= '0';
partial_product_10(87) <= '0';
partial_product_10(88) <= '0';
partial_product_10(89) <= '0';
partial_product_10(90) <= '0';
partial_product_10(91) <= '0';
partial_product_10(92) <= '0';
partial_product_10(93) <= '0';
partial_product_10(94) <= '0';
partial_product_10(95) <= '0';
partial_product_10(96) <= '0';
partial_product_10(97) <= '0';
partial_product_10(98) <= '0';
partial_product_10(99) <= '0';
partial_product_10(100) <= '0';
partial_product_10(101) <= '0';
partial_product_10(102) <= temp_mult_30(102);
partial_product_10(103) <= temp_mult_30(103);
partial_product_10(104) <= temp_mult_30(104);
partial_product_10(105) <= temp_mult_30(105);
partial_product_10(106) <= temp_mult_30(106);
partial_product_10(107) <= temp_mult_30(107);
partial_product_10(108) <= temp_mult_30(108);
partial_product_10(109) <= temp_mult_30(109);
partial_product_10(110) <= temp_mult_30(110);
partial_product_10(111) <= temp_mult_30(111);
partial_product_10(112) <= temp_mult_30(112);
partial_product_10(113) <= temp_mult_30(113);
partial_product_10(114) <= temp_mult_30(114);
partial_product_10(115) <= temp_mult_30(115);
partial_product_10(116) <= temp_mult_30(116);
partial_product_10(117) <= temp_mult_30(117);
partial_product_10(118) <= temp_mult_30(118);
partial_product_10(119) <= temp_mult_30(119);
partial_product_10(120) <= temp_mult_30(120);
partial_product_10(121) <= temp_mult_30(121);
partial_product_10(122) <= temp_mult_30(122);
partial_product_10(123) <= temp_mult_30(123);
partial_product_10(124) <= temp_mult_30(124);
partial_product_10(125) <= temp_mult_30(125);
partial_product_10(126) <= temp_mult_30(126);
partial_product_10(127) <= temp_mult_30(127);
partial_product_10(128) <= temp_mult_30(128);
partial_product_10(129) <= temp_mult_30(129);
partial_product_10(130) <= temp_mult_30(130);
partial_product_10(131) <= temp_mult_30(131);
partial_product_10(132) <= temp_mult_30(132);
partial_product_10(133) <= temp_mult_30(133);
partial_product_10(134) <= temp_mult_30(134);
partial_product_10(135) <= temp_mult_30(135);
partial_product_10(136) <= temp_mult_30(136);
partial_product_10(137) <= temp_mult_30(137);
partial_product_10(138) <= temp_mult_30(138);
partial_product_10(139) <= temp_mult_30(139);
partial_product_10(140) <= temp_mult_30(140);
partial_product_10(141) <= temp_mult_30(141);
partial_product_10(142) <= temp_mult_30(142);
partial_product_10(143) <= temp_mult_36(143);
partial_product_10(144) <= temp_mult_36(144);
partial_product_10(145) <= temp_mult_36(145);
partial_product_10(146) <= temp_mult_36(146);
partial_product_10(147) <= temp_mult_36(147);
partial_product_10(148) <= temp_mult_36(148);
partial_product_10(149) <= temp_mult_36(149);
partial_product_10(150) <= temp_mult_36(150);
partial_product_10(151) <= temp_mult_36(151);
partial_product_10(152) <= temp_mult_36(152);
partial_product_10(153) <= temp_mult_36(153);
partial_product_10(154) <= temp_mult_36(154);
partial_product_10(155) <= temp_mult_36(155);
partial_product_10(156) <= temp_mult_36(156);
partial_product_10(157) <= temp_mult_36(157);
partial_product_10(158) <= temp_mult_36(158);
partial_product_10(159) <= temp_mult_36(159);
partial_product_10(160) <= temp_mult_36(160);
partial_product_10(161) <= temp_mult_36(161);
partial_product_10(162) <= temp_mult_36(162);
partial_product_10(163) <= temp_mult_36(163);
partial_product_10(164) <= temp_mult_36(164);
partial_product_10(165) <= temp_mult_36(165);
partial_product_10(166) <= temp_mult_36(166);
partial_product_10(167) <= temp_mult_36(167);
partial_product_10(168) <= temp_mult_36(168);
partial_product_10(169) <= temp_mult_36(169);
partial_product_10(170) <= temp_mult_36(170);
partial_product_10(171) <= temp_mult_36(171);
partial_product_10(172) <= temp_mult_36(172);
partial_product_10(173) <= temp_mult_36(173);
partial_product_10(174) <= temp_mult_36(174);
partial_product_10(175) <= temp_mult_36(175);
partial_product_10(176) <= temp_mult_36(176);
partial_product_10(177) <= temp_mult_36(177);
partial_product_10(178) <= temp_mult_36(178);
partial_product_10(179) <= temp_mult_36(179);
partial_product_10(180) <= temp_mult_36(180);
partial_product_10(181) <= temp_mult_36(181);
partial_product_10(182) <= temp_mult_36(182);
partial_product_10(183) <= temp_mult_36(183);
partial_product_10(184) <= temp_mult_96(184);
partial_product_10(185) <= temp_mult_96(185);
partial_product_10(186) <= temp_mult_96(186);
partial_product_10(187) <= temp_mult_96(187);
partial_product_10(188) <= temp_mult_96(188);
partial_product_10(189) <= temp_mult_96(189);
partial_product_10(190) <= temp_mult_96(190);
partial_product_10(191) <= temp_mult_96(191);
partial_product_10(192) <= temp_mult_96(192);
partial_product_10(193) <= temp_mult_96(193);
partial_product_10(194) <= temp_mult_96(194);
partial_product_10(195) <= temp_mult_96(195);
partial_product_10(196) <= temp_mult_96(196);
partial_product_10(197) <= temp_mult_96(197);
partial_product_10(198) <= temp_mult_96(198);
partial_product_10(199) <= temp_mult_96(199);
partial_product_10(200) <= temp_mult_96(200);
partial_product_10(201) <= temp_mult_96(201);
partial_product_10(202) <= temp_mult_96(202);
partial_product_10(203) <= temp_mult_96(203);
partial_product_10(204) <= temp_mult_96(204);
partial_product_10(205) <= temp_mult_96(205);
partial_product_10(206) <= temp_mult_96(206);
partial_product_10(207) <= temp_mult_96(207);
partial_product_10(208) <= temp_mult_96(208);
partial_product_10(209) <= temp_mult_96(209);
partial_product_10(210) <= temp_mult_96(210);
partial_product_10(211) <= temp_mult_96(211);
partial_product_10(212) <= temp_mult_96(212);
partial_product_10(213) <= temp_mult_96(213);
partial_product_10(214) <= temp_mult_96(214);
partial_product_10(215) <= temp_mult_96(215);
partial_product_10(216) <= temp_mult_96(216);
partial_product_10(217) <= temp_mult_96(217);
partial_product_10(218) <= temp_mult_96(218);
partial_product_10(219) <= temp_mult_96(219);
partial_product_10(220) <= temp_mult_96(220);
partial_product_10(221) <= temp_mult_96(221);
partial_product_10(222) <= temp_mult_96(222);
partial_product_10(223) <= temp_mult_96(223);
partial_product_10(224) <= temp_mult_96(224);
partial_product_10(225) <= temp_mult_105(225);
partial_product_10(226) <= temp_mult_105(226);
partial_product_10(227) <= temp_mult_105(227);
partial_product_10(228) <= temp_mult_105(228);
partial_product_10(229) <= temp_mult_105(229);
partial_product_10(230) <= temp_mult_105(230);
partial_product_10(231) <= temp_mult_105(231);
partial_product_10(232) <= temp_mult_105(232);
partial_product_10(233) <= temp_mult_105(233);
partial_product_10(234) <= temp_mult_105(234);
partial_product_10(235) <= temp_mult_105(235);
partial_product_10(236) <= temp_mult_105(236);
partial_product_10(237) <= temp_mult_105(237);
partial_product_10(238) <= temp_mult_105(238);
partial_product_10(239) <= temp_mult_105(239);
partial_product_10(240) <= temp_mult_105(240);
partial_product_10(241) <= temp_mult_105(241);
partial_product_10(242) <= temp_mult_105(242);
partial_product_10(243) <= temp_mult_105(243);
partial_product_10(244) <= temp_mult_105(244);
partial_product_10(245) <= temp_mult_105(245);
partial_product_10(246) <= temp_mult_105(246);
partial_product_10(247) <= temp_mult_105(247);
partial_product_10(248) <= temp_mult_105(248);
partial_product_10(249) <= temp_mult_105(249);
partial_product_10(250) <= temp_mult_105(250);
partial_product_10(251) <= temp_mult_105(251);
partial_product_10(252) <= temp_mult_105(252);
partial_product_10(253) <= temp_mult_105(253);
partial_product_10(254) <= temp_mult_105(254);
partial_product_10(255) <= temp_mult_105(255);
partial_product_10(256) <= temp_mult_105(256);
partial_product_10(257) <= temp_mult_105(257);
partial_product_10(258) <= temp_mult_105(258);
partial_product_10(259) <= temp_mult_105(259);
partial_product_10(260) <= temp_mult_105(260);
partial_product_10(261) <= temp_mult_105(261);
partial_product_10(262) <= temp_mult_105(262);
partial_product_10(263) <= temp_mult_105(263);
partial_product_10(264) <= temp_mult_105(264);
partial_product_10(265) <= temp_mult_105(265);
partial_product_10(266) <= temp_mult_114(266);
partial_product_10(267) <= temp_mult_114(267);
partial_product_10(268) <= temp_mult_114(268);
partial_product_10(269) <= temp_mult_114(269);
partial_product_10(270) <= temp_mult_114(270);
partial_product_10(271) <= temp_mult_114(271);
partial_product_10(272) <= temp_mult_114(272);
partial_product_10(273) <= temp_mult_114(273);
partial_product_10(274) <= temp_mult_114(274);
partial_product_10(275) <= temp_mult_114(275);
partial_product_10(276) <= temp_mult_114(276);
partial_product_10(277) <= temp_mult_114(277);
partial_product_10(278) <= temp_mult_114(278);
partial_product_10(279) <= temp_mult_114(279);
partial_product_10(280) <= temp_mult_114(280);
partial_product_10(281) <= temp_mult_114(281);
partial_product_10(282) <= temp_mult_114(282);
partial_product_10(283) <= temp_mult_114(283);
partial_product_10(284) <= temp_mult_114(284);
partial_product_10(285) <= temp_mult_114(285);
partial_product_10(286) <= temp_mult_114(286);
partial_product_10(287) <= temp_mult_114(287);
partial_product_10(288) <= temp_mult_114(288);
partial_product_10(289) <= temp_mult_114(289);
partial_product_10(290) <= temp_mult_114(290);
partial_product_10(291) <= temp_mult_114(291);
partial_product_10(292) <= temp_mult_114(292);
partial_product_10(293) <= temp_mult_114(293);
partial_product_10(294) <= temp_mult_114(294);
partial_product_10(295) <= temp_mult_114(295);
partial_product_10(296) <= temp_mult_114(296);
partial_product_10(297) <= temp_mult_114(297);
partial_product_10(298) <= temp_mult_114(298);
partial_product_10(299) <= temp_mult_114(299);
partial_product_10(300) <= temp_mult_114(300);
partial_product_10(301) <= temp_mult_114(301);
partial_product_10(302) <= temp_mult_114(302);
partial_product_10(303) <= temp_mult_114(303);
partial_product_10(304) <= temp_mult_114(304);
partial_product_10(305) <= temp_mult_114(305);
partial_product_10(306) <= temp_mult_114(306);
partial_product_10(307) <= temp_mult_135(307);
partial_product_10(308) <= temp_mult_135(308);
partial_product_10(309) <= temp_mult_135(309);
partial_product_10(310) <= temp_mult_135(310);
partial_product_10(311) <= temp_mult_135(311);
partial_product_10(312) <= temp_mult_135(312);
partial_product_10(313) <= temp_mult_135(313);
partial_product_10(314) <= temp_mult_135(314);
partial_product_10(315) <= temp_mult_135(315);
partial_product_10(316) <= temp_mult_135(316);
partial_product_10(317) <= temp_mult_135(317);
partial_product_10(318) <= temp_mult_135(318);
partial_product_10(319) <= temp_mult_135(319);
partial_product_10(320) <= temp_mult_135(320);
partial_product_10(321) <= temp_mult_135(321);
partial_product_10(322) <= temp_mult_135(322);
partial_product_10(323) <= temp_mult_135(323);
partial_product_10(324) <= temp_mult_135(324);
partial_product_10(325) <= temp_mult_135(325);
partial_product_10(326) <= temp_mult_135(326);
partial_product_10(327) <= temp_mult_135(327);
partial_product_10(328) <= temp_mult_135(328);
partial_product_10(329) <= temp_mult_135(329);
partial_product_10(330) <= temp_mult_135(330);
partial_product_10(331) <= temp_mult_135(331);
partial_product_10(332) <= temp_mult_135(332);
partial_product_10(333) <= temp_mult_135(333);
partial_product_10(334) <= temp_mult_135(334);
partial_product_10(335) <= temp_mult_135(335);
partial_product_10(336) <= temp_mult_135(336);
partial_product_10(337) <= temp_mult_135(337);
partial_product_10(338) <= temp_mult_135(338);
partial_product_10(339) <= temp_mult_135(339);
partial_product_10(340) <= temp_mult_135(340);
partial_product_10(341) <= temp_mult_135(341);
partial_product_10(342) <= temp_mult_135(342);
partial_product_10(343) <= temp_mult_135(343);
partial_product_10(344) <= temp_mult_135(344);
partial_product_10(345) <= temp_mult_135(345);
partial_product_10(346) <= temp_mult_135(346);
partial_product_10(347) <= temp_mult_135(347);
partial_product_10(348) <= '0';
partial_product_10(349) <= '0';
partial_product_10(350) <= '0';
partial_product_10(351) <= temp_mult_119(351);
partial_product_10(352) <= temp_mult_119(352);
partial_product_10(353) <= temp_mult_119(353);
partial_product_10(354) <= temp_mult_119(354);
partial_product_10(355) <= temp_mult_119(355);
partial_product_10(356) <= temp_mult_119(356);
partial_product_10(357) <= temp_mult_119(357);
partial_product_10(358) <= temp_mult_119(358);
partial_product_10(359) <= temp_mult_119(359);
partial_product_10(360) <= temp_mult_119(360);
partial_product_10(361) <= temp_mult_119(361);
partial_product_10(362) <= temp_mult_119(362);
partial_product_10(363) <= temp_mult_119(363);
partial_product_10(364) <= temp_mult_119(364);
partial_product_10(365) <= temp_mult_119(365);
partial_product_10(366) <= temp_mult_119(366);
partial_product_10(367) <= temp_mult_119(367);
partial_product_10(368) <= temp_mult_119(368);
partial_product_10(369) <= temp_mult_119(369);
partial_product_10(370) <= temp_mult_119(370);
partial_product_10(371) <= temp_mult_119(371);
partial_product_10(372) <= temp_mult_119(372);
partial_product_10(373) <= temp_mult_119(373);
partial_product_10(374) <= temp_mult_119(374);
partial_product_10(375) <= temp_mult_119(375);
partial_product_10(376) <= temp_mult_119(376);
partial_product_10(377) <= temp_mult_119(377);
partial_product_10(378) <= temp_mult_119(378);
partial_product_10(379) <= temp_mult_119(379);
partial_product_10(380) <= temp_mult_119(380);
partial_product_10(381) <= temp_mult_119(381);
partial_product_10(382) <= temp_mult_119(382);
partial_product_10(383) <= temp_mult_119(383);
partial_product_10(384) <= temp_mult_119(384);
partial_product_10(385) <= temp_mult_119(385);
partial_product_10(386) <= temp_mult_119(386);
partial_product_10(387) <= temp_mult_119(387);
partial_product_10(388) <= temp_mult_119(388);
partial_product_10(389) <= temp_mult_119(389);
partial_product_10(390) <= temp_mult_119(390);
partial_product_10(391) <= temp_mult_119(391);
partial_product_10(392) <= '0';
partial_product_10(393) <= '0';
partial_product_10(394) <= '0';
partial_product_10(395) <= '0';
partial_product_10(396) <= '0';
partial_product_10(397) <= '0';
partial_product_10(398) <= '0';
partial_product_10(399) <= '0';
partial_product_10(400) <= '0';
partial_product_10(401) <= '0';
partial_product_10(402) <= '0';
partial_product_10(403) <= '0';
partial_product_10(404) <= '0';
partial_product_10(405) <= '0';
partial_product_10(406) <= '0';
partial_product_10(407) <= '0';
partial_product_10(408) <= '0';
partial_product_10(409) <= '0';
partial_product_10(410) <= '0';
partial_product_10(411) <= '0';
partial_product_10(412) <= '0';
partial_product_10(413) <= '0';
partial_product_10(414) <= '0';
partial_product_10(415) <= '0';
partial_product_10(416) <= '0';
partial_product_10(417) <= '0';
partial_product_10(418) <= '0';
partial_product_10(419) <= '0';
partial_product_10(420) <= '0';
partial_product_10(421) <= '0';
partial_product_10(422) <= '0';
partial_product_10(423) <= '0';
partial_product_10(424) <= '0';
partial_product_10(425) <= '0';
partial_product_10(426) <= '0';
partial_product_10(427) <= '0';
partial_product_10(428) <= '0';
partial_product_10(429) <= '0';
partial_product_10(430) <= '0';
partial_product_10(431) <= '0';
partial_product_10(432) <= '0';
partial_product_10(433) <= '0';
partial_product_10(434) <= '0';
partial_product_10(435) <= '0';
partial_product_10(436) <= '0';
partial_product_10(437) <= '0';
partial_product_10(438) <= '0';
partial_product_10(439) <= '0';
partial_product_10(440) <= '0';
partial_product_10(441) <= '0';
partial_product_10(442) <= '0';
partial_product_10(443) <= '0';
partial_product_10(444) <= '0';
partial_product_10(445) <= '0';
partial_product_10(446) <= '0';
partial_product_10(447) <= '0';
partial_product_10(448) <= '0';
partial_product_10(449) <= '0';
partial_product_10(450) <= '0';
partial_product_10(451) <= '0';
partial_product_10(452) <= '0';
partial_product_10(453) <= '0';
partial_product_10(454) <= '0';
partial_product_10(455) <= '0';
partial_product_10(456) <= '0';
partial_product_10(457) <= '0';
partial_product_10(458) <= '0';
partial_product_10(459) <= '0';
partial_product_10(460) <= '0';
partial_product_10(461) <= '0';
partial_product_10(462) <= '0';
partial_product_10(463) <= '0';
partial_product_10(464) <= '0';
partial_product_10(465) <= '0';
partial_product_10(466) <= '0';
partial_product_10(467) <= '0';
partial_product_10(468) <= '0';
partial_product_10(469) <= '0';
partial_product_10(470) <= '0';
partial_product_10(471) <= '0';
partial_product_10(472) <= '0';
partial_product_10(473) <= '0';
partial_product_10(474) <= '0';
partial_product_10(475) <= '0';
partial_product_10(476) <= '0';
partial_product_10(477) <= '0';
partial_product_10(478) <= '0';
partial_product_10(479) <= '0';
partial_product_10(480) <= '0';
partial_product_10(481) <= '0';
partial_product_10(482) <= '0';
partial_product_10(483) <= '0';
partial_product_10(484) <= '0';
partial_product_10(485) <= '0';
partial_product_10(486) <= '0';
partial_product_10(487) <= '0';
partial_product_10(488) <= '0';
partial_product_10(489) <= '0';
partial_product_10(490) <= '0';
partial_product_10(491) <= '0';
partial_product_10(492) <= '0';
partial_product_10(493) <= '0';
partial_product_10(494) <= '0';
partial_product_10(495) <= '0';
partial_product_10(496) <= '0';
partial_product_10(497) <= '0';
partial_product_10(498) <= '0';
partial_product_10(499) <= '0';
partial_product_10(500) <= '0';
partial_product_10(501) <= '0';
partial_product_10(502) <= '0';
partial_product_10(503) <= '0';
partial_product_10(504) <= '0';
partial_product_10(505) <= '0';
partial_product_10(506) <= '0';
partial_product_10(507) <= '0';
partial_product_10(508) <= '0';
partial_product_10(509) <= '0';
partial_product_10(510) <= '0';
partial_product_10(511) <= '0';
partial_product_10(512) <= '0';
partial_product_11(0) <= '0';
partial_product_11(1) <= '0';
partial_product_11(2) <= '0';
partial_product_11(3) <= '0';
partial_product_11(4) <= '0';
partial_product_11(5) <= '0';
partial_product_11(6) <= '0';
partial_product_11(7) <= '0';
partial_product_11(8) <= '0';
partial_product_11(9) <= '0';
partial_product_11(10) <= '0';
partial_product_11(11) <= '0';
partial_product_11(12) <= '0';
partial_product_11(13) <= '0';
partial_product_11(14) <= '0';
partial_product_11(15) <= '0';
partial_product_11(16) <= '0';
partial_product_11(17) <= '0';
partial_product_11(18) <= '0';
partial_product_11(19) <= '0';
partial_product_11(20) <= '0';
partial_product_11(21) <= '0';
partial_product_11(22) <= '0';
partial_product_11(23) <= '0';
partial_product_11(24) <= '0';
partial_product_11(25) <= '0';
partial_product_11(26) <= '0';
partial_product_11(27) <= '0';
partial_product_11(28) <= '0';
partial_product_11(29) <= '0';
partial_product_11(30) <= '0';
partial_product_11(31) <= '0';
partial_product_11(32) <= '0';
partial_product_11(33) <= '0';
partial_product_11(34) <= '0';
partial_product_11(35) <= '0';
partial_product_11(36) <= '0';
partial_product_11(37) <= '0';
partial_product_11(38) <= '0';
partial_product_11(39) <= '0';
partial_product_11(40) <= '0';
partial_product_11(41) <= '0';
partial_product_11(42) <= '0';
partial_product_11(43) <= '0';
partial_product_11(44) <= '0';
partial_product_11(45) <= '0';
partial_product_11(46) <= '0';
partial_product_11(47) <= '0';
partial_product_11(48) <= '0';
partial_product_11(49) <= '0';
partial_product_11(50) <= '0';
partial_product_11(51) <= '0';
partial_product_11(52) <= '0';
partial_product_11(53) <= '0';
partial_product_11(54) <= '0';
partial_product_11(55) <= '0';
partial_product_11(56) <= '0';
partial_product_11(57) <= '0';
partial_product_11(58) <= '0';
partial_product_11(59) <= '0';
partial_product_11(60) <= '0';
partial_product_11(61) <= '0';
partial_product_11(62) <= '0';
partial_product_11(63) <= '0';
partial_product_11(64) <= '0';
partial_product_11(65) <= '0';
partial_product_11(66) <= '0';
partial_product_11(67) <= '0';
partial_product_11(68) <= '0';
partial_product_11(69) <= '0';
partial_product_11(70) <= '0';
partial_product_11(71) <= '0';
partial_product_11(72) <= '0';
partial_product_11(73) <= '0';
partial_product_11(74) <= '0';
partial_product_11(75) <= '0';
partial_product_11(76) <= '0';
partial_product_11(77) <= '0';
partial_product_11(78) <= '0';
partial_product_11(79) <= '0';
partial_product_11(80) <= '0';
partial_product_11(81) <= '0';
partial_product_11(82) <= '0';
partial_product_11(83) <= '0';
partial_product_11(84) <= '0';
partial_product_11(85) <= '0';
partial_product_11(86) <= '0';
partial_product_11(87) <= '0';
partial_product_11(88) <= '0';
partial_product_11(89) <= '0';
partial_product_11(90) <= '0';
partial_product_11(91) <= '0';
partial_product_11(92) <= '0';
partial_product_11(93) <= '0';
partial_product_11(94) <= '0';
partial_product_11(95) <= '0';
partial_product_11(96) <= '0';
partial_product_11(97) <= '0';
partial_product_11(98) <= '0';
partial_product_11(99) <= '0';
partial_product_11(100) <= '0';
partial_product_11(101) <= '0';
partial_product_11(102) <= '0';
partial_product_11(103) <= '0';
partial_product_11(104) <= '0';
partial_product_11(105) <= '0';
partial_product_11(106) <= '0';
partial_product_11(107) <= '0';
partial_product_11(108) <= '0';
partial_product_11(109) <= '0';
partial_product_11(110) <= '0';
partial_product_11(111) <= '0';
partial_product_11(112) <= '0';
partial_product_11(113) <= '0';
partial_product_11(114) <= '0';
partial_product_11(115) <= '0';
partial_product_11(116) <= '0';
partial_product_11(117) <= '0';
partial_product_11(118) <= '0';
partial_product_11(119) <= temp_mult_35(119);
partial_product_11(120) <= temp_mult_35(120);
partial_product_11(121) <= temp_mult_35(121);
partial_product_11(122) <= temp_mult_35(122);
partial_product_11(123) <= temp_mult_35(123);
partial_product_11(124) <= temp_mult_35(124);
partial_product_11(125) <= temp_mult_35(125);
partial_product_11(126) <= temp_mult_35(126);
partial_product_11(127) <= temp_mult_35(127);
partial_product_11(128) <= temp_mult_35(128);
partial_product_11(129) <= temp_mult_35(129);
partial_product_11(130) <= temp_mult_35(130);
partial_product_11(131) <= temp_mult_35(131);
partial_product_11(132) <= temp_mult_35(132);
partial_product_11(133) <= temp_mult_35(133);
partial_product_11(134) <= temp_mult_35(134);
partial_product_11(135) <= temp_mult_35(135);
partial_product_11(136) <= temp_mult_35(136);
partial_product_11(137) <= temp_mult_35(137);
partial_product_11(138) <= temp_mult_35(138);
partial_product_11(139) <= temp_mult_35(139);
partial_product_11(140) <= temp_mult_35(140);
partial_product_11(141) <= temp_mult_35(141);
partial_product_11(142) <= temp_mult_35(142);
partial_product_11(143) <= temp_mult_35(143);
partial_product_11(144) <= temp_mult_35(144);
partial_product_11(145) <= temp_mult_35(145);
partial_product_11(146) <= temp_mult_35(146);
partial_product_11(147) <= temp_mult_35(147);
partial_product_11(148) <= temp_mult_35(148);
partial_product_11(149) <= temp_mult_35(149);
partial_product_11(150) <= temp_mult_35(150);
partial_product_11(151) <= temp_mult_35(151);
partial_product_11(152) <= temp_mult_35(152);
partial_product_11(153) <= temp_mult_35(153);
partial_product_11(154) <= temp_mult_35(154);
partial_product_11(155) <= temp_mult_35(155);
partial_product_11(156) <= temp_mult_35(156);
partial_product_11(157) <= temp_mult_35(157);
partial_product_11(158) <= temp_mult_35(158);
partial_product_11(159) <= temp_mult_35(159);
partial_product_11(160) <= temp_mult_88(160);
partial_product_11(161) <= temp_mult_88(161);
partial_product_11(162) <= temp_mult_88(162);
partial_product_11(163) <= temp_mult_88(163);
partial_product_11(164) <= temp_mult_88(164);
partial_product_11(165) <= temp_mult_88(165);
partial_product_11(166) <= temp_mult_88(166);
partial_product_11(167) <= temp_mult_88(167);
partial_product_11(168) <= temp_mult_88(168);
partial_product_11(169) <= temp_mult_88(169);
partial_product_11(170) <= temp_mult_88(170);
partial_product_11(171) <= temp_mult_88(171);
partial_product_11(172) <= temp_mult_88(172);
partial_product_11(173) <= temp_mult_88(173);
partial_product_11(174) <= temp_mult_88(174);
partial_product_11(175) <= temp_mult_88(175);
partial_product_11(176) <= temp_mult_88(176);
partial_product_11(177) <= temp_mult_88(177);
partial_product_11(178) <= temp_mult_88(178);
partial_product_11(179) <= temp_mult_88(179);
partial_product_11(180) <= temp_mult_88(180);
partial_product_11(181) <= temp_mult_88(181);
partial_product_11(182) <= temp_mult_88(182);
partial_product_11(183) <= temp_mult_88(183);
partial_product_11(184) <= temp_mult_88(184);
partial_product_11(185) <= temp_mult_88(185);
partial_product_11(186) <= temp_mult_88(186);
partial_product_11(187) <= temp_mult_88(187);
partial_product_11(188) <= temp_mult_88(188);
partial_product_11(189) <= temp_mult_88(189);
partial_product_11(190) <= temp_mult_88(190);
partial_product_11(191) <= temp_mult_88(191);
partial_product_11(192) <= temp_mult_88(192);
partial_product_11(193) <= temp_mult_88(193);
partial_product_11(194) <= temp_mult_88(194);
partial_product_11(195) <= temp_mult_88(195);
partial_product_11(196) <= temp_mult_88(196);
partial_product_11(197) <= temp_mult_88(197);
partial_product_11(198) <= temp_mult_88(198);
partial_product_11(199) <= temp_mult_88(199);
partial_product_11(200) <= temp_mult_88(200);
partial_product_11(201) <= temp_mult_97(201);
partial_product_11(202) <= temp_mult_97(202);
partial_product_11(203) <= temp_mult_97(203);
partial_product_11(204) <= temp_mult_97(204);
partial_product_11(205) <= temp_mult_97(205);
partial_product_11(206) <= temp_mult_97(206);
partial_product_11(207) <= temp_mult_97(207);
partial_product_11(208) <= temp_mult_97(208);
partial_product_11(209) <= temp_mult_97(209);
partial_product_11(210) <= temp_mult_97(210);
partial_product_11(211) <= temp_mult_97(211);
partial_product_11(212) <= temp_mult_97(212);
partial_product_11(213) <= temp_mult_97(213);
partial_product_11(214) <= temp_mult_97(214);
partial_product_11(215) <= temp_mult_97(215);
partial_product_11(216) <= temp_mult_97(216);
partial_product_11(217) <= temp_mult_97(217);
partial_product_11(218) <= temp_mult_97(218);
partial_product_11(219) <= temp_mult_97(219);
partial_product_11(220) <= temp_mult_97(220);
partial_product_11(221) <= temp_mult_97(221);
partial_product_11(222) <= temp_mult_97(222);
partial_product_11(223) <= temp_mult_97(223);
partial_product_11(224) <= temp_mult_97(224);
partial_product_11(225) <= temp_mult_97(225);
partial_product_11(226) <= temp_mult_97(226);
partial_product_11(227) <= temp_mult_97(227);
partial_product_11(228) <= temp_mult_97(228);
partial_product_11(229) <= temp_mult_97(229);
partial_product_11(230) <= temp_mult_97(230);
partial_product_11(231) <= temp_mult_97(231);
partial_product_11(232) <= temp_mult_97(232);
partial_product_11(233) <= temp_mult_97(233);
partial_product_11(234) <= temp_mult_97(234);
partial_product_11(235) <= temp_mult_97(235);
partial_product_11(236) <= temp_mult_97(236);
partial_product_11(237) <= temp_mult_97(237);
partial_product_11(238) <= temp_mult_97(238);
partial_product_11(239) <= temp_mult_97(239);
partial_product_11(240) <= temp_mult_97(240);
partial_product_11(241) <= temp_mult_97(241);
partial_product_11(242) <= temp_mult_106(242);
partial_product_11(243) <= temp_mult_106(243);
partial_product_11(244) <= temp_mult_106(244);
partial_product_11(245) <= temp_mult_106(245);
partial_product_11(246) <= temp_mult_106(246);
partial_product_11(247) <= temp_mult_106(247);
partial_product_11(248) <= temp_mult_106(248);
partial_product_11(249) <= temp_mult_106(249);
partial_product_11(250) <= temp_mult_106(250);
partial_product_11(251) <= temp_mult_106(251);
partial_product_11(252) <= temp_mult_106(252);
partial_product_11(253) <= temp_mult_106(253);
partial_product_11(254) <= temp_mult_106(254);
partial_product_11(255) <= temp_mult_106(255);
partial_product_11(256) <= temp_mult_106(256);
partial_product_11(257) <= temp_mult_106(257);
partial_product_11(258) <= temp_mult_106(258);
partial_product_11(259) <= temp_mult_106(259);
partial_product_11(260) <= temp_mult_106(260);
partial_product_11(261) <= temp_mult_106(261);
partial_product_11(262) <= temp_mult_106(262);
partial_product_11(263) <= temp_mult_106(263);
partial_product_11(264) <= temp_mult_106(264);
partial_product_11(265) <= temp_mult_106(265);
partial_product_11(266) <= temp_mult_106(266);
partial_product_11(267) <= temp_mult_106(267);
partial_product_11(268) <= temp_mult_106(268);
partial_product_11(269) <= temp_mult_106(269);
partial_product_11(270) <= temp_mult_106(270);
partial_product_11(271) <= temp_mult_106(271);
partial_product_11(272) <= temp_mult_106(272);
partial_product_11(273) <= temp_mult_106(273);
partial_product_11(274) <= temp_mult_106(274);
partial_product_11(275) <= temp_mult_106(275);
partial_product_11(276) <= temp_mult_106(276);
partial_product_11(277) <= temp_mult_106(277);
partial_product_11(278) <= temp_mult_106(278);
partial_product_11(279) <= temp_mult_106(279);
partial_product_11(280) <= temp_mult_106(280);
partial_product_11(281) <= temp_mult_106(281);
partial_product_11(282) <= temp_mult_106(282);
partial_product_11(283) <= temp_mult_115(283);
partial_product_11(284) <= temp_mult_115(284);
partial_product_11(285) <= temp_mult_115(285);
partial_product_11(286) <= temp_mult_115(286);
partial_product_11(287) <= temp_mult_115(287);
partial_product_11(288) <= temp_mult_115(288);
partial_product_11(289) <= temp_mult_115(289);
partial_product_11(290) <= temp_mult_115(290);
partial_product_11(291) <= temp_mult_115(291);
partial_product_11(292) <= temp_mult_115(292);
partial_product_11(293) <= temp_mult_115(293);
partial_product_11(294) <= temp_mult_115(294);
partial_product_11(295) <= temp_mult_115(295);
partial_product_11(296) <= temp_mult_115(296);
partial_product_11(297) <= temp_mult_115(297);
partial_product_11(298) <= temp_mult_115(298);
partial_product_11(299) <= temp_mult_115(299);
partial_product_11(300) <= temp_mult_115(300);
partial_product_11(301) <= temp_mult_115(301);
partial_product_11(302) <= temp_mult_115(302);
partial_product_11(303) <= temp_mult_115(303);
partial_product_11(304) <= temp_mult_115(304);
partial_product_11(305) <= temp_mult_115(305);
partial_product_11(306) <= temp_mult_115(306);
partial_product_11(307) <= temp_mult_115(307);
partial_product_11(308) <= temp_mult_115(308);
partial_product_11(309) <= temp_mult_115(309);
partial_product_11(310) <= temp_mult_115(310);
partial_product_11(311) <= temp_mult_115(311);
partial_product_11(312) <= temp_mult_115(312);
partial_product_11(313) <= temp_mult_115(313);
partial_product_11(314) <= temp_mult_115(314);
partial_product_11(315) <= temp_mult_115(315);
partial_product_11(316) <= temp_mult_115(316);
partial_product_11(317) <= temp_mult_115(317);
partial_product_11(318) <= temp_mult_115(318);
partial_product_11(319) <= temp_mult_115(319);
partial_product_11(320) <= temp_mult_115(320);
partial_product_11(321) <= temp_mult_115(321);
partial_product_11(322) <= temp_mult_115(322);
partial_product_11(323) <= temp_mult_115(323);
partial_product_11(324) <= temp_mult_140(324);
partial_product_11(325) <= temp_mult_140(325);
partial_product_11(326) <= temp_mult_140(326);
partial_product_11(327) <= temp_mult_140(327);
partial_product_11(328) <= temp_mult_140(328);
partial_product_11(329) <= temp_mult_140(329);
partial_product_11(330) <= temp_mult_140(330);
partial_product_11(331) <= temp_mult_140(331);
partial_product_11(332) <= temp_mult_140(332);
partial_product_11(333) <= temp_mult_140(333);
partial_product_11(334) <= temp_mult_140(334);
partial_product_11(335) <= temp_mult_140(335);
partial_product_11(336) <= temp_mult_140(336);
partial_product_11(337) <= temp_mult_140(337);
partial_product_11(338) <= temp_mult_140(338);
partial_product_11(339) <= temp_mult_140(339);
partial_product_11(340) <= temp_mult_140(340);
partial_product_11(341) <= temp_mult_140(341);
partial_product_11(342) <= temp_mult_140(342);
partial_product_11(343) <= temp_mult_140(343);
partial_product_11(344) <= temp_mult_140(344);
partial_product_11(345) <= temp_mult_140(345);
partial_product_11(346) <= temp_mult_140(346);
partial_product_11(347) <= temp_mult_140(347);
partial_product_11(348) <= temp_mult_140(348);
partial_product_11(349) <= temp_mult_140(349);
partial_product_11(350) <= temp_mult_140(350);
partial_product_11(351) <= temp_mult_140(351);
partial_product_11(352) <= temp_mult_140(352);
partial_product_11(353) <= temp_mult_140(353);
partial_product_11(354) <= temp_mult_140(354);
partial_product_11(355) <= temp_mult_140(355);
partial_product_11(356) <= temp_mult_140(356);
partial_product_11(357) <= temp_mult_140(357);
partial_product_11(358) <= temp_mult_140(358);
partial_product_11(359) <= temp_mult_140(359);
partial_product_11(360) <= temp_mult_140(360);
partial_product_11(361) <= temp_mult_140(361);
partial_product_11(362) <= temp_mult_140(362);
partial_product_11(363) <= temp_mult_140(363);
partial_product_11(364) <= temp_mult_140(364);
partial_product_11(365) <= '0';
partial_product_11(366) <= '0';
partial_product_11(367) <= '0';
partial_product_11(368) <= '0';
partial_product_11(369) <= '0';
partial_product_11(370) <= '0';
partial_product_11(371) <= '0';
partial_product_11(372) <= '0';
partial_product_11(373) <= '0';
partial_product_11(374) <= '0';
partial_product_11(375) <= temp_mult_155(375);
partial_product_11(376) <= temp_mult_155(376);
partial_product_11(377) <= temp_mult_155(377);
partial_product_11(378) <= temp_mult_155(378);
partial_product_11(379) <= temp_mult_155(379);
partial_product_11(380) <= temp_mult_155(380);
partial_product_11(381) <= temp_mult_155(381);
partial_product_11(382) <= temp_mult_155(382);
partial_product_11(383) <= temp_mult_155(383);
partial_product_11(384) <= temp_mult_155(384);
partial_product_11(385) <= temp_mult_155(385);
partial_product_11(386) <= temp_mult_155(386);
partial_product_11(387) <= temp_mult_155(387);
partial_product_11(388) <= temp_mult_155(388);
partial_product_11(389) <= temp_mult_155(389);
partial_product_11(390) <= temp_mult_155(390);
partial_product_11(391) <= temp_mult_155(391);
partial_product_11(392) <= temp_mult_155(392);
partial_product_11(393) <= temp_mult_155(393);
partial_product_11(394) <= temp_mult_155(394);
partial_product_11(395) <= temp_mult_155(395);
partial_product_11(396) <= temp_mult_155(396);
partial_product_11(397) <= temp_mult_155(397);
partial_product_11(398) <= temp_mult_155(398);
partial_product_11(399) <= temp_mult_155(399);
partial_product_11(400) <= temp_mult_155(400);
partial_product_11(401) <= temp_mult_155(401);
partial_product_11(402) <= temp_mult_155(402);
partial_product_11(403) <= temp_mult_155(403);
partial_product_11(404) <= temp_mult_155(404);
partial_product_11(405) <= temp_mult_155(405);
partial_product_11(406) <= temp_mult_155(406);
partial_product_11(407) <= temp_mult_155(407);
partial_product_11(408) <= temp_mult_155(408);
partial_product_11(409) <= temp_mult_155(409);
partial_product_11(410) <= temp_mult_155(410);
partial_product_11(411) <= temp_mult_155(411);
partial_product_11(412) <= temp_mult_155(412);
partial_product_11(413) <= temp_mult_155(413);
partial_product_11(414) <= temp_mult_155(414);
partial_product_11(415) <= temp_mult_155(415);
partial_product_11(416) <= '0';
partial_product_11(417) <= '0';
partial_product_11(418) <= '0';
partial_product_11(419) <= '0';
partial_product_11(420) <= '0';
partial_product_11(421) <= '0';
partial_product_11(422) <= '0';
partial_product_11(423) <= '0';
partial_product_11(424) <= '0';
partial_product_11(425) <= '0';
partial_product_11(426) <= '0';
partial_product_11(427) <= '0';
partial_product_11(428) <= '0';
partial_product_11(429) <= '0';
partial_product_11(430) <= '0';
partial_product_11(431) <= '0';
partial_product_11(432) <= '0';
partial_product_11(433) <= '0';
partial_product_11(434) <= '0';
partial_product_11(435) <= '0';
partial_product_11(436) <= '0';
partial_product_11(437) <= '0';
partial_product_11(438) <= '0';
partial_product_11(439) <= '0';
partial_product_11(440) <= '0';
partial_product_11(441) <= '0';
partial_product_11(442) <= '0';
partial_product_11(443) <= '0';
partial_product_11(444) <= '0';
partial_product_11(445) <= '0';
partial_product_11(446) <= '0';
partial_product_11(447) <= '0';
partial_product_11(448) <= '0';
partial_product_11(449) <= '0';
partial_product_11(450) <= '0';
partial_product_11(451) <= '0';
partial_product_11(452) <= '0';
partial_product_11(453) <= '0';
partial_product_11(454) <= '0';
partial_product_11(455) <= '0';
partial_product_11(456) <= '0';
partial_product_11(457) <= '0';
partial_product_11(458) <= '0';
partial_product_11(459) <= '0';
partial_product_11(460) <= '0';
partial_product_11(461) <= '0';
partial_product_11(462) <= '0';
partial_product_11(463) <= '0';
partial_product_11(464) <= '0';
partial_product_11(465) <= '0';
partial_product_11(466) <= '0';
partial_product_11(467) <= '0';
partial_product_11(468) <= '0';
partial_product_11(469) <= '0';
partial_product_11(470) <= '0';
partial_product_11(471) <= '0';
partial_product_11(472) <= '0';
partial_product_11(473) <= '0';
partial_product_11(474) <= '0';
partial_product_11(475) <= '0';
partial_product_11(476) <= '0';
partial_product_11(477) <= '0';
partial_product_11(478) <= '0';
partial_product_11(479) <= '0';
partial_product_11(480) <= '0';
partial_product_11(481) <= '0';
partial_product_11(482) <= '0';
partial_product_11(483) <= '0';
partial_product_11(484) <= '0';
partial_product_11(485) <= '0';
partial_product_11(486) <= '0';
partial_product_11(487) <= '0';
partial_product_11(488) <= '0';
partial_product_11(489) <= '0';
partial_product_11(490) <= '0';
partial_product_11(491) <= '0';
partial_product_11(492) <= '0';
partial_product_11(493) <= '0';
partial_product_11(494) <= '0';
partial_product_11(495) <= '0';
partial_product_11(496) <= '0';
partial_product_11(497) <= '0';
partial_product_11(498) <= '0';
partial_product_11(499) <= '0';
partial_product_11(500) <= '0';
partial_product_11(501) <= '0';
partial_product_11(502) <= '0';
partial_product_11(503) <= '0';
partial_product_11(504) <= '0';
partial_product_11(505) <= '0';
partial_product_11(506) <= '0';
partial_product_11(507) <= '0';
partial_product_11(508) <= '0';
partial_product_11(509) <= '0';
partial_product_11(510) <= '0';
partial_product_11(511) <= '0';
partial_product_11(512) <= '0';
partial_product_12(0) <= '0';
partial_product_12(1) <= '0';
partial_product_12(2) <= '0';
partial_product_12(3) <= '0';
partial_product_12(4) <= '0';
partial_product_12(5) <= '0';
partial_product_12(6) <= '0';
partial_product_12(7) <= '0';
partial_product_12(8) <= '0';
partial_product_12(9) <= '0';
partial_product_12(10) <= '0';
partial_product_12(11) <= '0';
partial_product_12(12) <= '0';
partial_product_12(13) <= '0';
partial_product_12(14) <= '0';
partial_product_12(15) <= '0';
partial_product_12(16) <= '0';
partial_product_12(17) <= '0';
partial_product_12(18) <= '0';
partial_product_12(19) <= '0';
partial_product_12(20) <= '0';
partial_product_12(21) <= '0';
partial_product_12(22) <= '0';
partial_product_12(23) <= '0';
partial_product_12(24) <= '0';
partial_product_12(25) <= '0';
partial_product_12(26) <= '0';
partial_product_12(27) <= '0';
partial_product_12(28) <= '0';
partial_product_12(29) <= '0';
partial_product_12(30) <= '0';
partial_product_12(31) <= '0';
partial_product_12(32) <= '0';
partial_product_12(33) <= '0';
partial_product_12(34) <= '0';
partial_product_12(35) <= '0';
partial_product_12(36) <= '0';
partial_product_12(37) <= '0';
partial_product_12(38) <= '0';
partial_product_12(39) <= '0';
partial_product_12(40) <= '0';
partial_product_12(41) <= '0';
partial_product_12(42) <= '0';
partial_product_12(43) <= '0';
partial_product_12(44) <= '0';
partial_product_12(45) <= '0';
partial_product_12(46) <= '0';
partial_product_12(47) <= '0';
partial_product_12(48) <= '0';
partial_product_12(49) <= '0';
partial_product_12(50) <= '0';
partial_product_12(51) <= '0';
partial_product_12(52) <= '0';
partial_product_12(53) <= '0';
partial_product_12(54) <= '0';
partial_product_12(55) <= '0';
partial_product_12(56) <= '0';
partial_product_12(57) <= '0';
partial_product_12(58) <= '0';
partial_product_12(59) <= '0';
partial_product_12(60) <= '0';
partial_product_12(61) <= '0';
partial_product_12(62) <= '0';
partial_product_12(63) <= '0';
partial_product_12(64) <= '0';
partial_product_12(65) <= '0';
partial_product_12(66) <= '0';
partial_product_12(67) <= '0';
partial_product_12(68) <= '0';
partial_product_12(69) <= '0';
partial_product_12(70) <= '0';
partial_product_12(71) <= '0';
partial_product_12(72) <= '0';
partial_product_12(73) <= '0';
partial_product_12(74) <= '0';
partial_product_12(75) <= '0';
partial_product_12(76) <= '0';
partial_product_12(77) <= '0';
partial_product_12(78) <= '0';
partial_product_12(79) <= '0';
partial_product_12(80) <= '0';
partial_product_12(81) <= '0';
partial_product_12(82) <= '0';
partial_product_12(83) <= '0';
partial_product_12(84) <= '0';
partial_product_12(85) <= '0';
partial_product_12(86) <= '0';
partial_product_12(87) <= '0';
partial_product_12(88) <= '0';
partial_product_12(89) <= '0';
partial_product_12(90) <= '0';
partial_product_12(91) <= '0';
partial_product_12(92) <= '0';
partial_product_12(93) <= '0';
partial_product_12(94) <= '0';
partial_product_12(95) <= '0';
partial_product_12(96) <= '0';
partial_product_12(97) <= '0';
partial_product_12(98) <= '0';
partial_product_12(99) <= '0';
partial_product_12(100) <= '0';
partial_product_12(101) <= '0';
partial_product_12(102) <= '0';
partial_product_12(103) <= '0';
partial_product_12(104) <= '0';
partial_product_12(105) <= '0';
partial_product_12(106) <= '0';
partial_product_12(107) <= '0';
partial_product_12(108) <= '0';
partial_product_12(109) <= '0';
partial_product_12(110) <= '0';
partial_product_12(111) <= '0';
partial_product_12(112) <= '0';
partial_product_12(113) <= '0';
partial_product_12(114) <= '0';
partial_product_12(115) <= '0';
partial_product_12(116) <= '0';
partial_product_12(117) <= '0';
partial_product_12(118) <= '0';
partial_product_12(119) <= '0';
partial_product_12(120) <= temp_mult_40(120);
partial_product_12(121) <= temp_mult_40(121);
partial_product_12(122) <= temp_mult_40(122);
partial_product_12(123) <= temp_mult_40(123);
partial_product_12(124) <= temp_mult_40(124);
partial_product_12(125) <= temp_mult_40(125);
partial_product_12(126) <= temp_mult_40(126);
partial_product_12(127) <= temp_mult_40(127);
partial_product_12(128) <= temp_mult_40(128);
partial_product_12(129) <= temp_mult_40(129);
partial_product_12(130) <= temp_mult_40(130);
partial_product_12(131) <= temp_mult_40(131);
partial_product_12(132) <= temp_mult_40(132);
partial_product_12(133) <= temp_mult_40(133);
partial_product_12(134) <= temp_mult_40(134);
partial_product_12(135) <= temp_mult_40(135);
partial_product_12(136) <= temp_mult_40(136);
partial_product_12(137) <= temp_mult_40(137);
partial_product_12(138) <= temp_mult_40(138);
partial_product_12(139) <= temp_mult_40(139);
partial_product_12(140) <= temp_mult_40(140);
partial_product_12(141) <= temp_mult_40(141);
partial_product_12(142) <= temp_mult_40(142);
partial_product_12(143) <= temp_mult_40(143);
partial_product_12(144) <= temp_mult_40(144);
partial_product_12(145) <= temp_mult_40(145);
partial_product_12(146) <= temp_mult_40(146);
partial_product_12(147) <= temp_mult_40(147);
partial_product_12(148) <= temp_mult_40(148);
partial_product_12(149) <= temp_mult_40(149);
partial_product_12(150) <= temp_mult_40(150);
partial_product_12(151) <= temp_mult_40(151);
partial_product_12(152) <= temp_mult_40(152);
partial_product_12(153) <= temp_mult_40(153);
partial_product_12(154) <= temp_mult_40(154);
partial_product_12(155) <= temp_mult_40(155);
partial_product_12(156) <= temp_mult_40(156);
partial_product_12(157) <= temp_mult_40(157);
partial_product_12(158) <= temp_mult_40(158);
partial_product_12(159) <= temp_mult_40(159);
partial_product_12(160) <= temp_mult_40(160);
partial_product_12(161) <= temp_mult_49(161);
partial_product_12(162) <= temp_mult_49(162);
partial_product_12(163) <= temp_mult_49(163);
partial_product_12(164) <= temp_mult_49(164);
partial_product_12(165) <= temp_mult_49(165);
partial_product_12(166) <= temp_mult_49(166);
partial_product_12(167) <= temp_mult_49(167);
partial_product_12(168) <= temp_mult_49(168);
partial_product_12(169) <= temp_mult_49(169);
partial_product_12(170) <= temp_mult_49(170);
partial_product_12(171) <= temp_mult_49(171);
partial_product_12(172) <= temp_mult_49(172);
partial_product_12(173) <= temp_mult_49(173);
partial_product_12(174) <= temp_mult_49(174);
partial_product_12(175) <= temp_mult_49(175);
partial_product_12(176) <= temp_mult_49(176);
partial_product_12(177) <= temp_mult_49(177);
partial_product_12(178) <= temp_mult_49(178);
partial_product_12(179) <= temp_mult_49(179);
partial_product_12(180) <= temp_mult_49(180);
partial_product_12(181) <= temp_mult_49(181);
partial_product_12(182) <= temp_mult_49(182);
partial_product_12(183) <= temp_mult_49(183);
partial_product_12(184) <= temp_mult_49(184);
partial_product_12(185) <= temp_mult_49(185);
partial_product_12(186) <= temp_mult_49(186);
partial_product_12(187) <= temp_mult_49(187);
partial_product_12(188) <= temp_mult_49(188);
partial_product_12(189) <= temp_mult_49(189);
partial_product_12(190) <= temp_mult_49(190);
partial_product_12(191) <= temp_mult_49(191);
partial_product_12(192) <= temp_mult_49(192);
partial_product_12(193) <= temp_mult_49(193);
partial_product_12(194) <= temp_mult_49(194);
partial_product_12(195) <= temp_mult_49(195);
partial_product_12(196) <= temp_mult_49(196);
partial_product_12(197) <= temp_mult_49(197);
partial_product_12(198) <= temp_mult_49(198);
partial_product_12(199) <= temp_mult_49(199);
partial_product_12(200) <= temp_mult_49(200);
partial_product_12(201) <= temp_mult_49(201);
partial_product_12(202) <= temp_mult_58(202);
partial_product_12(203) <= temp_mult_58(203);
partial_product_12(204) <= temp_mult_58(204);
partial_product_12(205) <= temp_mult_58(205);
partial_product_12(206) <= temp_mult_58(206);
partial_product_12(207) <= temp_mult_58(207);
partial_product_12(208) <= temp_mult_58(208);
partial_product_12(209) <= temp_mult_58(209);
partial_product_12(210) <= temp_mult_58(210);
partial_product_12(211) <= temp_mult_58(211);
partial_product_12(212) <= temp_mult_58(212);
partial_product_12(213) <= temp_mult_58(213);
partial_product_12(214) <= temp_mult_58(214);
partial_product_12(215) <= temp_mult_58(215);
partial_product_12(216) <= temp_mult_58(216);
partial_product_12(217) <= temp_mult_58(217);
partial_product_12(218) <= temp_mult_58(218);
partial_product_12(219) <= temp_mult_58(219);
partial_product_12(220) <= temp_mult_58(220);
partial_product_12(221) <= temp_mult_58(221);
partial_product_12(222) <= temp_mult_58(222);
partial_product_12(223) <= temp_mult_58(223);
partial_product_12(224) <= temp_mult_58(224);
partial_product_12(225) <= temp_mult_58(225);
partial_product_12(226) <= temp_mult_58(226);
partial_product_12(227) <= temp_mult_58(227);
partial_product_12(228) <= temp_mult_58(228);
partial_product_12(229) <= temp_mult_58(229);
partial_product_12(230) <= temp_mult_58(230);
partial_product_12(231) <= temp_mult_58(231);
partial_product_12(232) <= temp_mult_58(232);
partial_product_12(233) <= temp_mult_58(233);
partial_product_12(234) <= temp_mult_58(234);
partial_product_12(235) <= temp_mult_58(235);
partial_product_12(236) <= temp_mult_58(236);
partial_product_12(237) <= temp_mult_58(237);
partial_product_12(238) <= temp_mult_58(238);
partial_product_12(239) <= temp_mult_58(239);
partial_product_12(240) <= temp_mult_58(240);
partial_product_12(241) <= temp_mult_58(241);
partial_product_12(242) <= temp_mult_58(242);
partial_product_12(243) <= temp_mult_67(243);
partial_product_12(244) <= temp_mult_67(244);
partial_product_12(245) <= temp_mult_67(245);
partial_product_12(246) <= temp_mult_67(246);
partial_product_12(247) <= temp_mult_67(247);
partial_product_12(248) <= temp_mult_67(248);
partial_product_12(249) <= temp_mult_67(249);
partial_product_12(250) <= temp_mult_67(250);
partial_product_12(251) <= temp_mult_67(251);
partial_product_12(252) <= temp_mult_67(252);
partial_product_12(253) <= temp_mult_67(253);
partial_product_12(254) <= temp_mult_67(254);
partial_product_12(255) <= temp_mult_67(255);
partial_product_12(256) <= temp_mult_67(256);
partial_product_12(257) <= temp_mult_67(257);
partial_product_12(258) <= temp_mult_67(258);
partial_product_12(259) <= temp_mult_67(259);
partial_product_12(260) <= temp_mult_67(260);
partial_product_12(261) <= temp_mult_67(261);
partial_product_12(262) <= temp_mult_67(262);
partial_product_12(263) <= temp_mult_67(263);
partial_product_12(264) <= temp_mult_67(264);
partial_product_12(265) <= temp_mult_67(265);
partial_product_12(266) <= temp_mult_67(266);
partial_product_12(267) <= temp_mult_67(267);
partial_product_12(268) <= temp_mult_67(268);
partial_product_12(269) <= temp_mult_67(269);
partial_product_12(270) <= temp_mult_67(270);
partial_product_12(271) <= temp_mult_67(271);
partial_product_12(272) <= temp_mult_67(272);
partial_product_12(273) <= temp_mult_67(273);
partial_product_12(274) <= temp_mult_67(274);
partial_product_12(275) <= temp_mult_67(275);
partial_product_12(276) <= temp_mult_67(276);
partial_product_12(277) <= temp_mult_67(277);
partial_product_12(278) <= temp_mult_67(278);
partial_product_12(279) <= temp_mult_67(279);
partial_product_12(280) <= temp_mult_67(280);
partial_product_12(281) <= temp_mult_67(281);
partial_product_12(282) <= temp_mult_67(282);
partial_product_12(283) <= temp_mult_67(283);
partial_product_12(284) <= temp_mult_76(284);
partial_product_12(285) <= temp_mult_76(285);
partial_product_12(286) <= temp_mult_76(286);
partial_product_12(287) <= temp_mult_76(287);
partial_product_12(288) <= temp_mult_76(288);
partial_product_12(289) <= temp_mult_76(289);
partial_product_12(290) <= temp_mult_76(290);
partial_product_12(291) <= temp_mult_76(291);
partial_product_12(292) <= temp_mult_76(292);
partial_product_12(293) <= temp_mult_76(293);
partial_product_12(294) <= temp_mult_76(294);
partial_product_12(295) <= temp_mult_76(295);
partial_product_12(296) <= temp_mult_76(296);
partial_product_12(297) <= temp_mult_76(297);
partial_product_12(298) <= temp_mult_76(298);
partial_product_12(299) <= temp_mult_76(299);
partial_product_12(300) <= temp_mult_76(300);
partial_product_12(301) <= temp_mult_76(301);
partial_product_12(302) <= temp_mult_76(302);
partial_product_12(303) <= temp_mult_76(303);
partial_product_12(304) <= temp_mult_76(304);
partial_product_12(305) <= temp_mult_76(305);
partial_product_12(306) <= temp_mult_76(306);
partial_product_12(307) <= temp_mult_76(307);
partial_product_12(308) <= temp_mult_76(308);
partial_product_12(309) <= temp_mult_76(309);
partial_product_12(310) <= temp_mult_76(310);
partial_product_12(311) <= temp_mult_76(311);
partial_product_12(312) <= temp_mult_76(312);
partial_product_12(313) <= temp_mult_76(313);
partial_product_12(314) <= temp_mult_76(314);
partial_product_12(315) <= temp_mult_76(315);
partial_product_12(316) <= temp_mult_76(316);
partial_product_12(317) <= temp_mult_76(317);
partial_product_12(318) <= temp_mult_76(318);
partial_product_12(319) <= temp_mult_76(319);
partial_product_12(320) <= temp_mult_76(320);
partial_product_12(321) <= temp_mult_76(321);
partial_product_12(322) <= temp_mult_76(322);
partial_product_12(323) <= temp_mult_76(323);
partial_product_12(324) <= temp_mult_76(324);
partial_product_12(325) <= '0';
partial_product_12(326) <= '0';
partial_product_12(327) <= temp_mult_111(327);
partial_product_12(328) <= temp_mult_111(328);
partial_product_12(329) <= temp_mult_111(329);
partial_product_12(330) <= temp_mult_111(330);
partial_product_12(331) <= temp_mult_111(331);
partial_product_12(332) <= temp_mult_111(332);
partial_product_12(333) <= temp_mult_111(333);
partial_product_12(334) <= temp_mult_111(334);
partial_product_12(335) <= temp_mult_111(335);
partial_product_12(336) <= temp_mult_111(336);
partial_product_12(337) <= temp_mult_111(337);
partial_product_12(338) <= temp_mult_111(338);
partial_product_12(339) <= temp_mult_111(339);
partial_product_12(340) <= temp_mult_111(340);
partial_product_12(341) <= temp_mult_111(341);
partial_product_12(342) <= temp_mult_111(342);
partial_product_12(343) <= temp_mult_111(343);
partial_product_12(344) <= temp_mult_111(344);
partial_product_12(345) <= temp_mult_111(345);
partial_product_12(346) <= temp_mult_111(346);
partial_product_12(347) <= temp_mult_111(347);
partial_product_12(348) <= temp_mult_111(348);
partial_product_12(349) <= temp_mult_111(349);
partial_product_12(350) <= temp_mult_111(350);
partial_product_12(351) <= temp_mult_111(351);
partial_product_12(352) <= temp_mult_111(352);
partial_product_12(353) <= temp_mult_111(353);
partial_product_12(354) <= temp_mult_111(354);
partial_product_12(355) <= temp_mult_111(355);
partial_product_12(356) <= temp_mult_111(356);
partial_product_12(357) <= temp_mult_111(357);
partial_product_12(358) <= temp_mult_111(358);
partial_product_12(359) <= temp_mult_111(359);
partial_product_12(360) <= temp_mult_111(360);
partial_product_12(361) <= temp_mult_111(361);
partial_product_12(362) <= temp_mult_111(362);
partial_product_12(363) <= temp_mult_111(363);
partial_product_12(364) <= temp_mult_111(364);
partial_product_12(365) <= temp_mult_111(365);
partial_product_12(366) <= temp_mult_111(366);
partial_product_12(367) <= temp_mult_111(367);
partial_product_12(368) <= '0';
partial_product_12(369) <= '0';
partial_product_12(370) <= '0';
partial_product_12(371) <= '0';
partial_product_12(372) <= '0';
partial_product_12(373) <= '0';
partial_product_12(374) <= '0';
partial_product_12(375) <= '0';
partial_product_12(376) <= '0';
partial_product_12(377) <= '0';
partial_product_12(378) <= '0';
partial_product_12(379) <= '0';
partial_product_12(380) <= '0';
partial_product_12(381) <= '0';
partial_product_12(382) <= '0';
partial_product_12(383) <= '0';
partial_product_12(384) <= '0';
partial_product_12(385) <= '0';
partial_product_12(386) <= '0';
partial_product_12(387) <= '0';
partial_product_12(388) <= '0';
partial_product_12(389) <= '0';
partial_product_12(390) <= '0';
partial_product_12(391) <= '0';
partial_product_12(392) <= '0';
partial_product_12(393) <= '0';
partial_product_12(394) <= '0';
partial_product_12(395) <= '0';
partial_product_12(396) <= '0';
partial_product_12(397) <= '0';
partial_product_12(398) <= '0';
partial_product_12(399) <= '0';
partial_product_12(400) <= '0';
partial_product_12(401) <= '0';
partial_product_12(402) <= '0';
partial_product_12(403) <= '0';
partial_product_12(404) <= '0';
partial_product_12(405) <= '0';
partial_product_12(406) <= '0';
partial_product_12(407) <= '0';
partial_product_12(408) <= '0';
partial_product_12(409) <= '0';
partial_product_12(410) <= '0';
partial_product_12(411) <= '0';
partial_product_12(412) <= '0';
partial_product_12(413) <= '0';
partial_product_12(414) <= '0';
partial_product_12(415) <= '0';
partial_product_12(416) <= '0';
partial_product_12(417) <= '0';
partial_product_12(418) <= '0';
partial_product_12(419) <= '0';
partial_product_12(420) <= '0';
partial_product_12(421) <= '0';
partial_product_12(422) <= '0';
partial_product_12(423) <= '0';
partial_product_12(424) <= '0';
partial_product_12(425) <= '0';
partial_product_12(426) <= '0';
partial_product_12(427) <= '0';
partial_product_12(428) <= '0';
partial_product_12(429) <= '0';
partial_product_12(430) <= '0';
partial_product_12(431) <= '0';
partial_product_12(432) <= '0';
partial_product_12(433) <= '0';
partial_product_12(434) <= '0';
partial_product_12(435) <= '0';
partial_product_12(436) <= '0';
partial_product_12(437) <= '0';
partial_product_12(438) <= '0';
partial_product_12(439) <= '0';
partial_product_12(440) <= '0';
partial_product_12(441) <= '0';
partial_product_12(442) <= '0';
partial_product_12(443) <= '0';
partial_product_12(444) <= '0';
partial_product_12(445) <= '0';
partial_product_12(446) <= '0';
partial_product_12(447) <= '0';
partial_product_12(448) <= '0';
partial_product_12(449) <= '0';
partial_product_12(450) <= '0';
partial_product_12(451) <= '0';
partial_product_12(452) <= '0';
partial_product_12(453) <= '0';
partial_product_12(454) <= '0';
partial_product_12(455) <= '0';
partial_product_12(456) <= '0';
partial_product_12(457) <= '0';
partial_product_12(458) <= '0';
partial_product_12(459) <= '0';
partial_product_12(460) <= '0';
partial_product_12(461) <= '0';
partial_product_12(462) <= '0';
partial_product_12(463) <= '0';
partial_product_12(464) <= '0';
partial_product_12(465) <= '0';
partial_product_12(466) <= '0';
partial_product_12(467) <= '0';
partial_product_12(468) <= '0';
partial_product_12(469) <= '0';
partial_product_12(470) <= '0';
partial_product_12(471) <= '0';
partial_product_12(472) <= '0';
partial_product_12(473) <= '0';
partial_product_12(474) <= '0';
partial_product_12(475) <= '0';
partial_product_12(476) <= '0';
partial_product_12(477) <= '0';
partial_product_12(478) <= '0';
partial_product_12(479) <= '0';
partial_product_12(480) <= '0';
partial_product_12(481) <= '0';
partial_product_12(482) <= '0';
partial_product_12(483) <= '0';
partial_product_12(484) <= '0';
partial_product_12(485) <= '0';
partial_product_12(486) <= '0';
partial_product_12(487) <= '0';
partial_product_12(488) <= '0';
partial_product_12(489) <= '0';
partial_product_12(490) <= '0';
partial_product_12(491) <= '0';
partial_product_12(492) <= '0';
partial_product_12(493) <= '0';
partial_product_12(494) <= '0';
partial_product_12(495) <= '0';
partial_product_12(496) <= '0';
partial_product_12(497) <= '0';
partial_product_12(498) <= '0';
partial_product_12(499) <= '0';
partial_product_12(500) <= '0';
partial_product_12(501) <= '0';
partial_product_12(502) <= '0';
partial_product_12(503) <= '0';
partial_product_12(504) <= '0';
partial_product_12(505) <= '0';
partial_product_12(506) <= '0';
partial_product_12(507) <= '0';
partial_product_12(508) <= '0';
partial_product_12(509) <= '0';
partial_product_12(510) <= '0';
partial_product_12(511) <= '0';
partial_product_12(512) <= '0';
partial_product_13(0) <= '0';
partial_product_13(1) <= '0';
partial_product_13(2) <= '0';
partial_product_13(3) <= '0';
partial_product_13(4) <= '0';
partial_product_13(5) <= '0';
partial_product_13(6) <= '0';
partial_product_13(7) <= '0';
partial_product_13(8) <= '0';
partial_product_13(9) <= '0';
partial_product_13(10) <= '0';
partial_product_13(11) <= '0';
partial_product_13(12) <= '0';
partial_product_13(13) <= '0';
partial_product_13(14) <= '0';
partial_product_13(15) <= '0';
partial_product_13(16) <= '0';
partial_product_13(17) <= '0';
partial_product_13(18) <= '0';
partial_product_13(19) <= '0';
partial_product_13(20) <= '0';
partial_product_13(21) <= '0';
partial_product_13(22) <= '0';
partial_product_13(23) <= '0';
partial_product_13(24) <= '0';
partial_product_13(25) <= '0';
partial_product_13(26) <= '0';
partial_product_13(27) <= '0';
partial_product_13(28) <= '0';
partial_product_13(29) <= '0';
partial_product_13(30) <= '0';
partial_product_13(31) <= '0';
partial_product_13(32) <= '0';
partial_product_13(33) <= '0';
partial_product_13(34) <= '0';
partial_product_13(35) <= '0';
partial_product_13(36) <= '0';
partial_product_13(37) <= '0';
partial_product_13(38) <= '0';
partial_product_13(39) <= '0';
partial_product_13(40) <= '0';
partial_product_13(41) <= '0';
partial_product_13(42) <= '0';
partial_product_13(43) <= '0';
partial_product_13(44) <= '0';
partial_product_13(45) <= '0';
partial_product_13(46) <= '0';
partial_product_13(47) <= '0';
partial_product_13(48) <= '0';
partial_product_13(49) <= '0';
partial_product_13(50) <= '0';
partial_product_13(51) <= '0';
partial_product_13(52) <= '0';
partial_product_13(53) <= '0';
partial_product_13(54) <= '0';
partial_product_13(55) <= '0';
partial_product_13(56) <= '0';
partial_product_13(57) <= '0';
partial_product_13(58) <= '0';
partial_product_13(59) <= '0';
partial_product_13(60) <= '0';
partial_product_13(61) <= '0';
partial_product_13(62) <= '0';
partial_product_13(63) <= '0';
partial_product_13(64) <= '0';
partial_product_13(65) <= '0';
partial_product_13(66) <= '0';
partial_product_13(67) <= '0';
partial_product_13(68) <= '0';
partial_product_13(69) <= '0';
partial_product_13(70) <= '0';
partial_product_13(71) <= '0';
partial_product_13(72) <= '0';
partial_product_13(73) <= '0';
partial_product_13(74) <= '0';
partial_product_13(75) <= '0';
partial_product_13(76) <= '0';
partial_product_13(77) <= '0';
partial_product_13(78) <= '0';
partial_product_13(79) <= '0';
partial_product_13(80) <= '0';
partial_product_13(81) <= '0';
partial_product_13(82) <= '0';
partial_product_13(83) <= '0';
partial_product_13(84) <= '0';
partial_product_13(85) <= '0';
partial_product_13(86) <= '0';
partial_product_13(87) <= '0';
partial_product_13(88) <= '0';
partial_product_13(89) <= '0';
partial_product_13(90) <= '0';
partial_product_13(91) <= '0';
partial_product_13(92) <= '0';
partial_product_13(93) <= '0';
partial_product_13(94) <= '0';
partial_product_13(95) <= '0';
partial_product_13(96) <= '0';
partial_product_13(97) <= '0';
partial_product_13(98) <= '0';
partial_product_13(99) <= '0';
partial_product_13(100) <= '0';
partial_product_13(101) <= '0';
partial_product_13(102) <= '0';
partial_product_13(103) <= '0';
partial_product_13(104) <= '0';
partial_product_13(105) <= '0';
partial_product_13(106) <= '0';
partial_product_13(107) <= '0';
partial_product_13(108) <= '0';
partial_product_13(109) <= '0';
partial_product_13(110) <= '0';
partial_product_13(111) <= '0';
partial_product_13(112) <= '0';
partial_product_13(113) <= '0';
partial_product_13(114) <= '0';
partial_product_13(115) <= '0';
partial_product_13(116) <= '0';
partial_product_13(117) <= '0';
partial_product_13(118) <= '0';
partial_product_13(119) <= '0';
partial_product_13(120) <= '0';
partial_product_13(121) <= '0';
partial_product_13(122) <= '0';
partial_product_13(123) <= '0';
partial_product_13(124) <= '0';
partial_product_13(125) <= '0';
partial_product_13(126) <= '0';
partial_product_13(127) <= '0';
partial_product_13(128) <= '0';
partial_product_13(129) <= '0';
partial_product_13(130) <= '0';
partial_product_13(131) <= '0';
partial_product_13(132) <= '0';
partial_product_13(133) <= '0';
partial_product_13(134) <= '0';
partial_product_13(135) <= '0';
partial_product_13(136) <= temp_mult_80(136);
partial_product_13(137) <= temp_mult_80(137);
partial_product_13(138) <= temp_mult_80(138);
partial_product_13(139) <= temp_mult_80(139);
partial_product_13(140) <= temp_mult_80(140);
partial_product_13(141) <= temp_mult_80(141);
partial_product_13(142) <= temp_mult_80(142);
partial_product_13(143) <= temp_mult_80(143);
partial_product_13(144) <= temp_mult_80(144);
partial_product_13(145) <= temp_mult_80(145);
partial_product_13(146) <= temp_mult_80(146);
partial_product_13(147) <= temp_mult_80(147);
partial_product_13(148) <= temp_mult_80(148);
partial_product_13(149) <= temp_mult_80(149);
partial_product_13(150) <= temp_mult_80(150);
partial_product_13(151) <= temp_mult_80(151);
partial_product_13(152) <= temp_mult_80(152);
partial_product_13(153) <= temp_mult_80(153);
partial_product_13(154) <= temp_mult_80(154);
partial_product_13(155) <= temp_mult_80(155);
partial_product_13(156) <= temp_mult_80(156);
partial_product_13(157) <= temp_mult_80(157);
partial_product_13(158) <= temp_mult_80(158);
partial_product_13(159) <= temp_mult_80(159);
partial_product_13(160) <= temp_mult_80(160);
partial_product_13(161) <= temp_mult_80(161);
partial_product_13(162) <= temp_mult_80(162);
partial_product_13(163) <= temp_mult_80(163);
partial_product_13(164) <= temp_mult_80(164);
partial_product_13(165) <= temp_mult_80(165);
partial_product_13(166) <= temp_mult_80(166);
partial_product_13(167) <= temp_mult_80(167);
partial_product_13(168) <= temp_mult_80(168);
partial_product_13(169) <= temp_mult_80(169);
partial_product_13(170) <= temp_mult_80(170);
partial_product_13(171) <= temp_mult_80(171);
partial_product_13(172) <= temp_mult_80(172);
partial_product_13(173) <= temp_mult_80(173);
partial_product_13(174) <= temp_mult_80(174);
partial_product_13(175) <= temp_mult_80(175);
partial_product_13(176) <= temp_mult_80(176);
partial_product_13(177) <= temp_mult_89(177);
partial_product_13(178) <= temp_mult_89(178);
partial_product_13(179) <= temp_mult_89(179);
partial_product_13(180) <= temp_mult_89(180);
partial_product_13(181) <= temp_mult_89(181);
partial_product_13(182) <= temp_mult_89(182);
partial_product_13(183) <= temp_mult_89(183);
partial_product_13(184) <= temp_mult_89(184);
partial_product_13(185) <= temp_mult_89(185);
partial_product_13(186) <= temp_mult_89(186);
partial_product_13(187) <= temp_mult_89(187);
partial_product_13(188) <= temp_mult_89(188);
partial_product_13(189) <= temp_mult_89(189);
partial_product_13(190) <= temp_mult_89(190);
partial_product_13(191) <= temp_mult_89(191);
partial_product_13(192) <= temp_mult_89(192);
partial_product_13(193) <= temp_mult_89(193);
partial_product_13(194) <= temp_mult_89(194);
partial_product_13(195) <= temp_mult_89(195);
partial_product_13(196) <= temp_mult_89(196);
partial_product_13(197) <= temp_mult_89(197);
partial_product_13(198) <= temp_mult_89(198);
partial_product_13(199) <= temp_mult_89(199);
partial_product_13(200) <= temp_mult_89(200);
partial_product_13(201) <= temp_mult_89(201);
partial_product_13(202) <= temp_mult_89(202);
partial_product_13(203) <= temp_mult_89(203);
partial_product_13(204) <= temp_mult_89(204);
partial_product_13(205) <= temp_mult_89(205);
partial_product_13(206) <= temp_mult_89(206);
partial_product_13(207) <= temp_mult_89(207);
partial_product_13(208) <= temp_mult_89(208);
partial_product_13(209) <= temp_mult_89(209);
partial_product_13(210) <= temp_mult_89(210);
partial_product_13(211) <= temp_mult_89(211);
partial_product_13(212) <= temp_mult_89(212);
partial_product_13(213) <= temp_mult_89(213);
partial_product_13(214) <= temp_mult_89(214);
partial_product_13(215) <= temp_mult_89(215);
partial_product_13(216) <= temp_mult_89(216);
partial_product_13(217) <= temp_mult_89(217);
partial_product_13(218) <= temp_mult_98(218);
partial_product_13(219) <= temp_mult_98(219);
partial_product_13(220) <= temp_mult_98(220);
partial_product_13(221) <= temp_mult_98(221);
partial_product_13(222) <= temp_mult_98(222);
partial_product_13(223) <= temp_mult_98(223);
partial_product_13(224) <= temp_mult_98(224);
partial_product_13(225) <= temp_mult_98(225);
partial_product_13(226) <= temp_mult_98(226);
partial_product_13(227) <= temp_mult_98(227);
partial_product_13(228) <= temp_mult_98(228);
partial_product_13(229) <= temp_mult_98(229);
partial_product_13(230) <= temp_mult_98(230);
partial_product_13(231) <= temp_mult_98(231);
partial_product_13(232) <= temp_mult_98(232);
partial_product_13(233) <= temp_mult_98(233);
partial_product_13(234) <= temp_mult_98(234);
partial_product_13(235) <= temp_mult_98(235);
partial_product_13(236) <= temp_mult_98(236);
partial_product_13(237) <= temp_mult_98(237);
partial_product_13(238) <= temp_mult_98(238);
partial_product_13(239) <= temp_mult_98(239);
partial_product_13(240) <= temp_mult_98(240);
partial_product_13(241) <= temp_mult_98(241);
partial_product_13(242) <= temp_mult_98(242);
partial_product_13(243) <= temp_mult_98(243);
partial_product_13(244) <= temp_mult_98(244);
partial_product_13(245) <= temp_mult_98(245);
partial_product_13(246) <= temp_mult_98(246);
partial_product_13(247) <= temp_mult_98(247);
partial_product_13(248) <= temp_mult_98(248);
partial_product_13(249) <= temp_mult_98(249);
partial_product_13(250) <= temp_mult_98(250);
partial_product_13(251) <= temp_mult_98(251);
partial_product_13(252) <= temp_mult_98(252);
partial_product_13(253) <= temp_mult_98(253);
partial_product_13(254) <= temp_mult_98(254);
partial_product_13(255) <= temp_mult_98(255);
partial_product_13(256) <= temp_mult_98(256);
partial_product_13(257) <= temp_mult_98(257);
partial_product_13(258) <= temp_mult_98(258);
partial_product_13(259) <= temp_mult_107(259);
partial_product_13(260) <= temp_mult_107(260);
partial_product_13(261) <= temp_mult_107(261);
partial_product_13(262) <= temp_mult_107(262);
partial_product_13(263) <= temp_mult_107(263);
partial_product_13(264) <= temp_mult_107(264);
partial_product_13(265) <= temp_mult_107(265);
partial_product_13(266) <= temp_mult_107(266);
partial_product_13(267) <= temp_mult_107(267);
partial_product_13(268) <= temp_mult_107(268);
partial_product_13(269) <= temp_mult_107(269);
partial_product_13(270) <= temp_mult_107(270);
partial_product_13(271) <= temp_mult_107(271);
partial_product_13(272) <= temp_mult_107(272);
partial_product_13(273) <= temp_mult_107(273);
partial_product_13(274) <= temp_mult_107(274);
partial_product_13(275) <= temp_mult_107(275);
partial_product_13(276) <= temp_mult_107(276);
partial_product_13(277) <= temp_mult_107(277);
partial_product_13(278) <= temp_mult_107(278);
partial_product_13(279) <= temp_mult_107(279);
partial_product_13(280) <= temp_mult_107(280);
partial_product_13(281) <= temp_mult_107(281);
partial_product_13(282) <= temp_mult_107(282);
partial_product_13(283) <= temp_mult_107(283);
partial_product_13(284) <= temp_mult_107(284);
partial_product_13(285) <= temp_mult_107(285);
partial_product_13(286) <= temp_mult_107(286);
partial_product_13(287) <= temp_mult_107(287);
partial_product_13(288) <= temp_mult_107(288);
partial_product_13(289) <= temp_mult_107(289);
partial_product_13(290) <= temp_mult_107(290);
partial_product_13(291) <= temp_mult_107(291);
partial_product_13(292) <= temp_mult_107(292);
partial_product_13(293) <= temp_mult_107(293);
partial_product_13(294) <= temp_mult_107(294);
partial_product_13(295) <= temp_mult_107(295);
partial_product_13(296) <= temp_mult_107(296);
partial_product_13(297) <= temp_mult_107(297);
partial_product_13(298) <= temp_mult_107(298);
partial_product_13(299) <= temp_mult_107(299);
partial_product_13(300) <= temp_mult_116(300);
partial_product_13(301) <= temp_mult_116(301);
partial_product_13(302) <= temp_mult_116(302);
partial_product_13(303) <= temp_mult_116(303);
partial_product_13(304) <= temp_mult_116(304);
partial_product_13(305) <= temp_mult_116(305);
partial_product_13(306) <= temp_mult_116(306);
partial_product_13(307) <= temp_mult_116(307);
partial_product_13(308) <= temp_mult_116(308);
partial_product_13(309) <= temp_mult_116(309);
partial_product_13(310) <= temp_mult_116(310);
partial_product_13(311) <= temp_mult_116(311);
partial_product_13(312) <= temp_mult_116(312);
partial_product_13(313) <= temp_mult_116(313);
partial_product_13(314) <= temp_mult_116(314);
partial_product_13(315) <= temp_mult_116(315);
partial_product_13(316) <= temp_mult_116(316);
partial_product_13(317) <= temp_mult_116(317);
partial_product_13(318) <= temp_mult_116(318);
partial_product_13(319) <= temp_mult_116(319);
partial_product_13(320) <= temp_mult_116(320);
partial_product_13(321) <= temp_mult_116(321);
partial_product_13(322) <= temp_mult_116(322);
partial_product_13(323) <= temp_mult_116(323);
partial_product_13(324) <= temp_mult_116(324);
partial_product_13(325) <= temp_mult_116(325);
partial_product_13(326) <= temp_mult_116(326);
partial_product_13(327) <= temp_mult_116(327);
partial_product_13(328) <= temp_mult_116(328);
partial_product_13(329) <= temp_mult_116(329);
partial_product_13(330) <= temp_mult_116(330);
partial_product_13(331) <= temp_mult_116(331);
partial_product_13(332) <= temp_mult_116(332);
partial_product_13(333) <= temp_mult_116(333);
partial_product_13(334) <= temp_mult_116(334);
partial_product_13(335) <= temp_mult_116(335);
partial_product_13(336) <= temp_mult_116(336);
partial_product_13(337) <= temp_mult_116(337);
partial_product_13(338) <= temp_mult_116(338);
partial_product_13(339) <= temp_mult_116(339);
partial_product_13(340) <= temp_mult_116(340);
partial_product_13(341) <= temp_mult_145(341);
partial_product_13(342) <= temp_mult_145(342);
partial_product_13(343) <= temp_mult_145(343);
partial_product_13(344) <= temp_mult_145(344);
partial_product_13(345) <= temp_mult_145(345);
partial_product_13(346) <= temp_mult_145(346);
partial_product_13(347) <= temp_mult_145(347);
partial_product_13(348) <= temp_mult_145(348);
partial_product_13(349) <= temp_mult_145(349);
partial_product_13(350) <= temp_mult_145(350);
partial_product_13(351) <= temp_mult_145(351);
partial_product_13(352) <= temp_mult_145(352);
partial_product_13(353) <= temp_mult_145(353);
partial_product_13(354) <= temp_mult_145(354);
partial_product_13(355) <= temp_mult_145(355);
partial_product_13(356) <= temp_mult_145(356);
partial_product_13(357) <= temp_mult_145(357);
partial_product_13(358) <= temp_mult_145(358);
partial_product_13(359) <= temp_mult_145(359);
partial_product_13(360) <= temp_mult_145(360);
partial_product_13(361) <= temp_mult_145(361);
partial_product_13(362) <= temp_mult_145(362);
partial_product_13(363) <= temp_mult_145(363);
partial_product_13(364) <= temp_mult_145(364);
partial_product_13(365) <= temp_mult_145(365);
partial_product_13(366) <= temp_mult_145(366);
partial_product_13(367) <= temp_mult_145(367);
partial_product_13(368) <= temp_mult_145(368);
partial_product_13(369) <= temp_mult_145(369);
partial_product_13(370) <= temp_mult_145(370);
partial_product_13(371) <= temp_mult_145(371);
partial_product_13(372) <= temp_mult_145(372);
partial_product_13(373) <= temp_mult_145(373);
partial_product_13(374) <= temp_mult_145(374);
partial_product_13(375) <= temp_mult_145(375);
partial_product_13(376) <= temp_mult_145(376);
partial_product_13(377) <= temp_mult_145(377);
partial_product_13(378) <= temp_mult_145(378);
partial_product_13(379) <= temp_mult_145(379);
partial_product_13(380) <= temp_mult_145(380);
partial_product_13(381) <= temp_mult_145(381);
partial_product_13(382) <= '0';
partial_product_13(383) <= '0';
partial_product_13(384) <= '0';
partial_product_13(385) <= '0';
partial_product_13(386) <= '0';
partial_product_13(387) <= '0';
partial_product_13(388) <= '0';
partial_product_13(389) <= '0';
partial_product_13(390) <= '0';
partial_product_13(391) <= '0';
partial_product_13(392) <= '0';
partial_product_13(393) <= '0';
partial_product_13(394) <= '0';
partial_product_13(395) <= '0';
partial_product_13(396) <= '0';
partial_product_13(397) <= '0';
partial_product_13(398) <= '0';
partial_product_13(399) <= '0';
partial_product_13(400) <= '0';
partial_product_13(401) <= '0';
partial_product_13(402) <= '0';
partial_product_13(403) <= '0';
partial_product_13(404) <= '0';
partial_product_13(405) <= '0';
partial_product_13(406) <= '0';
partial_product_13(407) <= '0';
partial_product_13(408) <= '0';
partial_product_13(409) <= '0';
partial_product_13(410) <= '0';
partial_product_13(411) <= '0';
partial_product_13(412) <= '0';
partial_product_13(413) <= '0';
partial_product_13(414) <= '0';
partial_product_13(415) <= '0';
partial_product_13(416) <= '0';
partial_product_13(417) <= '0';
partial_product_13(418) <= '0';
partial_product_13(419) <= '0';
partial_product_13(420) <= '0';
partial_product_13(421) <= '0';
partial_product_13(422) <= '0';
partial_product_13(423) <= '0';
partial_product_13(424) <= '0';
partial_product_13(425) <= '0';
partial_product_13(426) <= '0';
partial_product_13(427) <= '0';
partial_product_13(428) <= '0';
partial_product_13(429) <= '0';
partial_product_13(430) <= '0';
partial_product_13(431) <= '0';
partial_product_13(432) <= '0';
partial_product_13(433) <= '0';
partial_product_13(434) <= '0';
partial_product_13(435) <= '0';
partial_product_13(436) <= '0';
partial_product_13(437) <= '0';
partial_product_13(438) <= '0';
partial_product_13(439) <= '0';
partial_product_13(440) <= '0';
partial_product_13(441) <= '0';
partial_product_13(442) <= '0';
partial_product_13(443) <= '0';
partial_product_13(444) <= '0';
partial_product_13(445) <= '0';
partial_product_13(446) <= '0';
partial_product_13(447) <= '0';
partial_product_13(448) <= '0';
partial_product_13(449) <= '0';
partial_product_13(450) <= '0';
partial_product_13(451) <= '0';
partial_product_13(452) <= '0';
partial_product_13(453) <= '0';
partial_product_13(454) <= '0';
partial_product_13(455) <= '0';
partial_product_13(456) <= '0';
partial_product_13(457) <= '0';
partial_product_13(458) <= '0';
partial_product_13(459) <= '0';
partial_product_13(460) <= '0';
partial_product_13(461) <= '0';
partial_product_13(462) <= '0';
partial_product_13(463) <= '0';
partial_product_13(464) <= '0';
partial_product_13(465) <= '0';
partial_product_13(466) <= '0';
partial_product_13(467) <= '0';
partial_product_13(468) <= '0';
partial_product_13(469) <= '0';
partial_product_13(470) <= '0';
partial_product_13(471) <= '0';
partial_product_13(472) <= '0';
partial_product_13(473) <= '0';
partial_product_13(474) <= '0';
partial_product_13(475) <= '0';
partial_product_13(476) <= '0';
partial_product_13(477) <= '0';
partial_product_13(478) <= '0';
partial_product_13(479) <= '0';
partial_product_13(480) <= '0';
partial_product_13(481) <= '0';
partial_product_13(482) <= '0';
partial_product_13(483) <= '0';
partial_product_13(484) <= '0';
partial_product_13(485) <= '0';
partial_product_13(486) <= '0';
partial_product_13(487) <= '0';
partial_product_13(488) <= '0';
partial_product_13(489) <= '0';
partial_product_13(490) <= '0';
partial_product_13(491) <= '0';
partial_product_13(492) <= '0';
partial_product_13(493) <= '0';
partial_product_13(494) <= '0';
partial_product_13(495) <= '0';
partial_product_13(496) <= '0';
partial_product_13(497) <= '0';
partial_product_13(498) <= '0';
partial_product_13(499) <= '0';
partial_product_13(500) <= '0';
partial_product_13(501) <= '0';
partial_product_13(502) <= '0';
partial_product_13(503) <= '0';
partial_product_13(504) <= '0';
partial_product_13(505) <= '0';
partial_product_13(506) <= '0';
partial_product_13(507) <= '0';
partial_product_13(508) <= '0';
partial_product_13(509) <= '0';
partial_product_13(510) <= '0';
partial_product_13(511) <= '0';
partial_product_13(512) <= '0';
partial_product_14(0) <= '0';
partial_product_14(1) <= '0';
partial_product_14(2) <= '0';
partial_product_14(3) <= '0';
partial_product_14(4) <= '0';
partial_product_14(5) <= '0';
partial_product_14(6) <= '0';
partial_product_14(7) <= '0';
partial_product_14(8) <= '0';
partial_product_14(9) <= '0';
partial_product_14(10) <= '0';
partial_product_14(11) <= '0';
partial_product_14(12) <= '0';
partial_product_14(13) <= '0';
partial_product_14(14) <= '0';
partial_product_14(15) <= '0';
partial_product_14(16) <= '0';
partial_product_14(17) <= '0';
partial_product_14(18) <= '0';
partial_product_14(19) <= '0';
partial_product_14(20) <= '0';
partial_product_14(21) <= '0';
partial_product_14(22) <= '0';
partial_product_14(23) <= '0';
partial_product_14(24) <= '0';
partial_product_14(25) <= '0';
partial_product_14(26) <= '0';
partial_product_14(27) <= '0';
partial_product_14(28) <= '0';
partial_product_14(29) <= '0';
partial_product_14(30) <= '0';
partial_product_14(31) <= '0';
partial_product_14(32) <= '0';
partial_product_14(33) <= '0';
partial_product_14(34) <= '0';
partial_product_14(35) <= '0';
partial_product_14(36) <= '0';
partial_product_14(37) <= '0';
partial_product_14(38) <= '0';
partial_product_14(39) <= '0';
partial_product_14(40) <= '0';
partial_product_14(41) <= '0';
partial_product_14(42) <= '0';
partial_product_14(43) <= '0';
partial_product_14(44) <= '0';
partial_product_14(45) <= '0';
partial_product_14(46) <= '0';
partial_product_14(47) <= '0';
partial_product_14(48) <= '0';
partial_product_14(49) <= '0';
partial_product_14(50) <= '0';
partial_product_14(51) <= '0';
partial_product_14(52) <= '0';
partial_product_14(53) <= '0';
partial_product_14(54) <= '0';
partial_product_14(55) <= '0';
partial_product_14(56) <= '0';
partial_product_14(57) <= '0';
partial_product_14(58) <= '0';
partial_product_14(59) <= '0';
partial_product_14(60) <= '0';
partial_product_14(61) <= '0';
partial_product_14(62) <= '0';
partial_product_14(63) <= '0';
partial_product_14(64) <= '0';
partial_product_14(65) <= '0';
partial_product_14(66) <= '0';
partial_product_14(67) <= '0';
partial_product_14(68) <= '0';
partial_product_14(69) <= '0';
partial_product_14(70) <= '0';
partial_product_14(71) <= '0';
partial_product_14(72) <= '0';
partial_product_14(73) <= '0';
partial_product_14(74) <= '0';
partial_product_14(75) <= '0';
partial_product_14(76) <= '0';
partial_product_14(77) <= '0';
partial_product_14(78) <= '0';
partial_product_14(79) <= '0';
partial_product_14(80) <= '0';
partial_product_14(81) <= '0';
partial_product_14(82) <= '0';
partial_product_14(83) <= '0';
partial_product_14(84) <= '0';
partial_product_14(85) <= '0';
partial_product_14(86) <= '0';
partial_product_14(87) <= '0';
partial_product_14(88) <= '0';
partial_product_14(89) <= '0';
partial_product_14(90) <= '0';
partial_product_14(91) <= '0';
partial_product_14(92) <= '0';
partial_product_14(93) <= '0';
partial_product_14(94) <= '0';
partial_product_14(95) <= '0';
partial_product_14(96) <= '0';
partial_product_14(97) <= '0';
partial_product_14(98) <= '0';
partial_product_14(99) <= '0';
partial_product_14(100) <= '0';
partial_product_14(101) <= '0';
partial_product_14(102) <= '0';
partial_product_14(103) <= '0';
partial_product_14(104) <= '0';
partial_product_14(105) <= '0';
partial_product_14(106) <= '0';
partial_product_14(107) <= '0';
partial_product_14(108) <= '0';
partial_product_14(109) <= '0';
partial_product_14(110) <= '0';
partial_product_14(111) <= '0';
partial_product_14(112) <= '0';
partial_product_14(113) <= '0';
partial_product_14(114) <= '0';
partial_product_14(115) <= '0';
partial_product_14(116) <= '0';
partial_product_14(117) <= '0';
partial_product_14(118) <= '0';
partial_product_14(119) <= '0';
partial_product_14(120) <= '0';
partial_product_14(121) <= '0';
partial_product_14(122) <= '0';
partial_product_14(123) <= '0';
partial_product_14(124) <= '0';
partial_product_14(125) <= '0';
partial_product_14(126) <= '0';
partial_product_14(127) <= '0';
partial_product_14(128) <= '0';
partial_product_14(129) <= '0';
partial_product_14(130) <= '0';
partial_product_14(131) <= '0';
partial_product_14(132) <= '0';
partial_product_14(133) <= '0';
partial_product_14(134) <= '0';
partial_product_14(135) <= '0';
partial_product_14(136) <= '0';
partial_product_14(137) <= '0';
partial_product_14(138) <= '0';
partial_product_14(139) <= '0';
partial_product_14(140) <= '0';
partial_product_14(141) <= '0';
partial_product_14(142) <= '0';
partial_product_14(143) <= '0';
partial_product_14(144) <= temp_mult_48(144);
partial_product_14(145) <= temp_mult_48(145);
partial_product_14(146) <= temp_mult_48(146);
partial_product_14(147) <= temp_mult_48(147);
partial_product_14(148) <= temp_mult_48(148);
partial_product_14(149) <= temp_mult_48(149);
partial_product_14(150) <= temp_mult_48(150);
partial_product_14(151) <= temp_mult_48(151);
partial_product_14(152) <= temp_mult_48(152);
partial_product_14(153) <= temp_mult_48(153);
partial_product_14(154) <= temp_mult_48(154);
partial_product_14(155) <= temp_mult_48(155);
partial_product_14(156) <= temp_mult_48(156);
partial_product_14(157) <= temp_mult_48(157);
partial_product_14(158) <= temp_mult_48(158);
partial_product_14(159) <= temp_mult_48(159);
partial_product_14(160) <= temp_mult_48(160);
partial_product_14(161) <= temp_mult_48(161);
partial_product_14(162) <= temp_mult_48(162);
partial_product_14(163) <= temp_mult_48(163);
partial_product_14(164) <= temp_mult_48(164);
partial_product_14(165) <= temp_mult_48(165);
partial_product_14(166) <= temp_mult_48(166);
partial_product_14(167) <= temp_mult_48(167);
partial_product_14(168) <= temp_mult_48(168);
partial_product_14(169) <= temp_mult_48(169);
partial_product_14(170) <= temp_mult_48(170);
partial_product_14(171) <= temp_mult_48(171);
partial_product_14(172) <= temp_mult_48(172);
partial_product_14(173) <= temp_mult_48(173);
partial_product_14(174) <= temp_mult_48(174);
partial_product_14(175) <= temp_mult_48(175);
partial_product_14(176) <= temp_mult_48(176);
partial_product_14(177) <= temp_mult_48(177);
partial_product_14(178) <= temp_mult_48(178);
partial_product_14(179) <= temp_mult_48(179);
partial_product_14(180) <= temp_mult_48(180);
partial_product_14(181) <= temp_mult_48(181);
partial_product_14(182) <= temp_mult_48(182);
partial_product_14(183) <= temp_mult_48(183);
partial_product_14(184) <= temp_mult_48(184);
partial_product_14(185) <= temp_mult_57(185);
partial_product_14(186) <= temp_mult_57(186);
partial_product_14(187) <= temp_mult_57(187);
partial_product_14(188) <= temp_mult_57(188);
partial_product_14(189) <= temp_mult_57(189);
partial_product_14(190) <= temp_mult_57(190);
partial_product_14(191) <= temp_mult_57(191);
partial_product_14(192) <= temp_mult_57(192);
partial_product_14(193) <= temp_mult_57(193);
partial_product_14(194) <= temp_mult_57(194);
partial_product_14(195) <= temp_mult_57(195);
partial_product_14(196) <= temp_mult_57(196);
partial_product_14(197) <= temp_mult_57(197);
partial_product_14(198) <= temp_mult_57(198);
partial_product_14(199) <= temp_mult_57(199);
partial_product_14(200) <= temp_mult_57(200);
partial_product_14(201) <= temp_mult_57(201);
partial_product_14(202) <= temp_mult_57(202);
partial_product_14(203) <= temp_mult_57(203);
partial_product_14(204) <= temp_mult_57(204);
partial_product_14(205) <= temp_mult_57(205);
partial_product_14(206) <= temp_mult_57(206);
partial_product_14(207) <= temp_mult_57(207);
partial_product_14(208) <= temp_mult_57(208);
partial_product_14(209) <= temp_mult_57(209);
partial_product_14(210) <= temp_mult_57(210);
partial_product_14(211) <= temp_mult_57(211);
partial_product_14(212) <= temp_mult_57(212);
partial_product_14(213) <= temp_mult_57(213);
partial_product_14(214) <= temp_mult_57(214);
partial_product_14(215) <= temp_mult_57(215);
partial_product_14(216) <= temp_mult_57(216);
partial_product_14(217) <= temp_mult_57(217);
partial_product_14(218) <= temp_mult_57(218);
partial_product_14(219) <= temp_mult_57(219);
partial_product_14(220) <= temp_mult_57(220);
partial_product_14(221) <= temp_mult_57(221);
partial_product_14(222) <= temp_mult_57(222);
partial_product_14(223) <= temp_mult_57(223);
partial_product_14(224) <= temp_mult_57(224);
partial_product_14(225) <= temp_mult_57(225);
partial_product_14(226) <= temp_mult_66(226);
partial_product_14(227) <= temp_mult_66(227);
partial_product_14(228) <= temp_mult_66(228);
partial_product_14(229) <= temp_mult_66(229);
partial_product_14(230) <= temp_mult_66(230);
partial_product_14(231) <= temp_mult_66(231);
partial_product_14(232) <= temp_mult_66(232);
partial_product_14(233) <= temp_mult_66(233);
partial_product_14(234) <= temp_mult_66(234);
partial_product_14(235) <= temp_mult_66(235);
partial_product_14(236) <= temp_mult_66(236);
partial_product_14(237) <= temp_mult_66(237);
partial_product_14(238) <= temp_mult_66(238);
partial_product_14(239) <= temp_mult_66(239);
partial_product_14(240) <= temp_mult_66(240);
partial_product_14(241) <= temp_mult_66(241);
partial_product_14(242) <= temp_mult_66(242);
partial_product_14(243) <= temp_mult_66(243);
partial_product_14(244) <= temp_mult_66(244);
partial_product_14(245) <= temp_mult_66(245);
partial_product_14(246) <= temp_mult_66(246);
partial_product_14(247) <= temp_mult_66(247);
partial_product_14(248) <= temp_mult_66(248);
partial_product_14(249) <= temp_mult_66(249);
partial_product_14(250) <= temp_mult_66(250);
partial_product_14(251) <= temp_mult_66(251);
partial_product_14(252) <= temp_mult_66(252);
partial_product_14(253) <= temp_mult_66(253);
partial_product_14(254) <= temp_mult_66(254);
partial_product_14(255) <= temp_mult_66(255);
partial_product_14(256) <= temp_mult_66(256);
partial_product_14(257) <= temp_mult_66(257);
partial_product_14(258) <= temp_mult_66(258);
partial_product_14(259) <= temp_mult_66(259);
partial_product_14(260) <= temp_mult_66(260);
partial_product_14(261) <= temp_mult_66(261);
partial_product_14(262) <= temp_mult_66(262);
partial_product_14(263) <= temp_mult_66(263);
partial_product_14(264) <= temp_mult_66(264);
partial_product_14(265) <= temp_mult_66(265);
partial_product_14(266) <= temp_mult_66(266);
partial_product_14(267) <= temp_mult_75(267);
partial_product_14(268) <= temp_mult_75(268);
partial_product_14(269) <= temp_mult_75(269);
partial_product_14(270) <= temp_mult_75(270);
partial_product_14(271) <= temp_mult_75(271);
partial_product_14(272) <= temp_mult_75(272);
partial_product_14(273) <= temp_mult_75(273);
partial_product_14(274) <= temp_mult_75(274);
partial_product_14(275) <= temp_mult_75(275);
partial_product_14(276) <= temp_mult_75(276);
partial_product_14(277) <= temp_mult_75(277);
partial_product_14(278) <= temp_mult_75(278);
partial_product_14(279) <= temp_mult_75(279);
partial_product_14(280) <= temp_mult_75(280);
partial_product_14(281) <= temp_mult_75(281);
partial_product_14(282) <= temp_mult_75(282);
partial_product_14(283) <= temp_mult_75(283);
partial_product_14(284) <= temp_mult_75(284);
partial_product_14(285) <= temp_mult_75(285);
partial_product_14(286) <= temp_mult_75(286);
partial_product_14(287) <= temp_mult_75(287);
partial_product_14(288) <= temp_mult_75(288);
partial_product_14(289) <= temp_mult_75(289);
partial_product_14(290) <= temp_mult_75(290);
partial_product_14(291) <= temp_mult_75(291);
partial_product_14(292) <= temp_mult_75(292);
partial_product_14(293) <= temp_mult_75(293);
partial_product_14(294) <= temp_mult_75(294);
partial_product_14(295) <= temp_mult_75(295);
partial_product_14(296) <= temp_mult_75(296);
partial_product_14(297) <= temp_mult_75(297);
partial_product_14(298) <= temp_mult_75(298);
partial_product_14(299) <= temp_mult_75(299);
partial_product_14(300) <= temp_mult_75(300);
partial_product_14(301) <= temp_mult_75(301);
partial_product_14(302) <= temp_mult_75(302);
partial_product_14(303) <= temp_mult_75(303);
partial_product_14(304) <= temp_mult_75(304);
partial_product_14(305) <= temp_mult_75(305);
partial_product_14(306) <= temp_mult_75(306);
partial_product_14(307) <= temp_mult_75(307);
partial_product_14(308) <= '0';
partial_product_14(309) <= '0';
partial_product_14(310) <= temp_mult_110(310);
partial_product_14(311) <= temp_mult_110(311);
partial_product_14(312) <= temp_mult_110(312);
partial_product_14(313) <= temp_mult_110(313);
partial_product_14(314) <= temp_mult_110(314);
partial_product_14(315) <= temp_mult_110(315);
partial_product_14(316) <= temp_mult_110(316);
partial_product_14(317) <= temp_mult_110(317);
partial_product_14(318) <= temp_mult_110(318);
partial_product_14(319) <= temp_mult_110(319);
partial_product_14(320) <= temp_mult_110(320);
partial_product_14(321) <= temp_mult_110(321);
partial_product_14(322) <= temp_mult_110(322);
partial_product_14(323) <= temp_mult_110(323);
partial_product_14(324) <= temp_mult_110(324);
partial_product_14(325) <= temp_mult_110(325);
partial_product_14(326) <= temp_mult_110(326);
partial_product_14(327) <= temp_mult_110(327);
partial_product_14(328) <= temp_mult_110(328);
partial_product_14(329) <= temp_mult_110(329);
partial_product_14(330) <= temp_mult_110(330);
partial_product_14(331) <= temp_mult_110(331);
partial_product_14(332) <= temp_mult_110(332);
partial_product_14(333) <= temp_mult_110(333);
partial_product_14(334) <= temp_mult_110(334);
partial_product_14(335) <= temp_mult_110(335);
partial_product_14(336) <= temp_mult_110(336);
partial_product_14(337) <= temp_mult_110(337);
partial_product_14(338) <= temp_mult_110(338);
partial_product_14(339) <= temp_mult_110(339);
partial_product_14(340) <= temp_mult_110(340);
partial_product_14(341) <= temp_mult_110(341);
partial_product_14(342) <= temp_mult_110(342);
partial_product_14(343) <= temp_mult_110(343);
partial_product_14(344) <= temp_mult_110(344);
partial_product_14(345) <= temp_mult_110(345);
partial_product_14(346) <= temp_mult_110(346);
partial_product_14(347) <= temp_mult_110(347);
partial_product_14(348) <= temp_mult_110(348);
partial_product_14(349) <= temp_mult_110(349);
partial_product_14(350) <= temp_mult_110(350);
partial_product_14(351) <= '0';
partial_product_14(352) <= '0';
partial_product_14(353) <= '0';
partial_product_14(354) <= '0';
partial_product_14(355) <= '0';
partial_product_14(356) <= '0';
partial_product_14(357) <= '0';
partial_product_14(358) <= temp_mult_150(358);
partial_product_14(359) <= temp_mult_150(359);
partial_product_14(360) <= temp_mult_150(360);
partial_product_14(361) <= temp_mult_150(361);
partial_product_14(362) <= temp_mult_150(362);
partial_product_14(363) <= temp_mult_150(363);
partial_product_14(364) <= temp_mult_150(364);
partial_product_14(365) <= temp_mult_150(365);
partial_product_14(366) <= temp_mult_150(366);
partial_product_14(367) <= temp_mult_150(367);
partial_product_14(368) <= temp_mult_150(368);
partial_product_14(369) <= temp_mult_150(369);
partial_product_14(370) <= temp_mult_150(370);
partial_product_14(371) <= temp_mult_150(371);
partial_product_14(372) <= temp_mult_150(372);
partial_product_14(373) <= temp_mult_150(373);
partial_product_14(374) <= temp_mult_150(374);
partial_product_14(375) <= temp_mult_150(375);
partial_product_14(376) <= temp_mult_150(376);
partial_product_14(377) <= temp_mult_150(377);
partial_product_14(378) <= temp_mult_150(378);
partial_product_14(379) <= temp_mult_150(379);
partial_product_14(380) <= temp_mult_150(380);
partial_product_14(381) <= temp_mult_150(381);
partial_product_14(382) <= temp_mult_150(382);
partial_product_14(383) <= temp_mult_150(383);
partial_product_14(384) <= temp_mult_150(384);
partial_product_14(385) <= temp_mult_150(385);
partial_product_14(386) <= temp_mult_150(386);
partial_product_14(387) <= temp_mult_150(387);
partial_product_14(388) <= temp_mult_150(388);
partial_product_14(389) <= temp_mult_150(389);
partial_product_14(390) <= temp_mult_150(390);
partial_product_14(391) <= temp_mult_150(391);
partial_product_14(392) <= temp_mult_150(392);
partial_product_14(393) <= temp_mult_150(393);
partial_product_14(394) <= temp_mult_150(394);
partial_product_14(395) <= temp_mult_150(395);
partial_product_14(396) <= temp_mult_150(396);
partial_product_14(397) <= temp_mult_150(397);
partial_product_14(398) <= temp_mult_150(398);
partial_product_14(399) <= '0';
partial_product_14(400) <= '0';
partial_product_14(401) <= '0';
partial_product_14(402) <= '0';
partial_product_14(403) <= '0';
partial_product_14(404) <= '0';
partial_product_14(405) <= '0';
partial_product_14(406) <= '0';
partial_product_14(407) <= '0';
partial_product_14(408) <= '0';
partial_product_14(409) <= '0';
partial_product_14(410) <= '0';
partial_product_14(411) <= '0';
partial_product_14(412) <= '0';
partial_product_14(413) <= '0';
partial_product_14(414) <= '0';
partial_product_14(415) <= '0';
partial_product_14(416) <= '0';
partial_product_14(417) <= '0';
partial_product_14(418) <= '0';
partial_product_14(419) <= '0';
partial_product_14(420) <= '0';
partial_product_14(421) <= '0';
partial_product_14(422) <= '0';
partial_product_14(423) <= '0';
partial_product_14(424) <= '0';
partial_product_14(425) <= '0';
partial_product_14(426) <= '0';
partial_product_14(427) <= '0';
partial_product_14(428) <= '0';
partial_product_14(429) <= '0';
partial_product_14(430) <= '0';
partial_product_14(431) <= '0';
partial_product_14(432) <= '0';
partial_product_14(433) <= '0';
partial_product_14(434) <= '0';
partial_product_14(435) <= '0';
partial_product_14(436) <= '0';
partial_product_14(437) <= '0';
partial_product_14(438) <= '0';
partial_product_14(439) <= '0';
partial_product_14(440) <= '0';
partial_product_14(441) <= '0';
partial_product_14(442) <= '0';
partial_product_14(443) <= '0';
partial_product_14(444) <= '0';
partial_product_14(445) <= '0';
partial_product_14(446) <= '0';
partial_product_14(447) <= '0';
partial_product_14(448) <= '0';
partial_product_14(449) <= '0';
partial_product_14(450) <= '0';
partial_product_14(451) <= '0';
partial_product_14(452) <= '0';
partial_product_14(453) <= '0';
partial_product_14(454) <= '0';
partial_product_14(455) <= '0';
partial_product_14(456) <= '0';
partial_product_14(457) <= '0';
partial_product_14(458) <= '0';
partial_product_14(459) <= '0';
partial_product_14(460) <= '0';
partial_product_14(461) <= '0';
partial_product_14(462) <= '0';
partial_product_14(463) <= '0';
partial_product_14(464) <= '0';
partial_product_14(465) <= '0';
partial_product_14(466) <= '0';
partial_product_14(467) <= '0';
partial_product_14(468) <= '0';
partial_product_14(469) <= '0';
partial_product_14(470) <= '0';
partial_product_14(471) <= '0';
partial_product_14(472) <= '0';
partial_product_14(473) <= '0';
partial_product_14(474) <= '0';
partial_product_14(475) <= '0';
partial_product_14(476) <= '0';
partial_product_14(477) <= '0';
partial_product_14(478) <= '0';
partial_product_14(479) <= '0';
partial_product_14(480) <= '0';
partial_product_14(481) <= '0';
partial_product_14(482) <= '0';
partial_product_14(483) <= '0';
partial_product_14(484) <= '0';
partial_product_14(485) <= '0';
partial_product_14(486) <= '0';
partial_product_14(487) <= '0';
partial_product_14(488) <= '0';
partial_product_14(489) <= '0';
partial_product_14(490) <= '0';
partial_product_14(491) <= '0';
partial_product_14(492) <= '0';
partial_product_14(493) <= '0';
partial_product_14(494) <= '0';
partial_product_14(495) <= '0';
partial_product_14(496) <= '0';
partial_product_14(497) <= '0';
partial_product_14(498) <= '0';
partial_product_14(499) <= '0';
partial_product_14(500) <= '0';
partial_product_14(501) <= '0';
partial_product_14(502) <= '0';
partial_product_14(503) <= '0';
partial_product_14(504) <= '0';
partial_product_14(505) <= '0';
partial_product_14(506) <= '0';
partial_product_14(507) <= '0';
partial_product_14(508) <= '0';
partial_product_14(509) <= '0';
partial_product_14(510) <= '0';
partial_product_14(511) <= '0';
partial_product_14(512) <= '0';
partial_product_15(0) <= '0';
partial_product_15(1) <= '0';
partial_product_15(2) <= '0';
partial_product_15(3) <= '0';
partial_product_15(4) <= '0';
partial_product_15(5) <= '0';
partial_product_15(6) <= '0';
partial_product_15(7) <= '0';
partial_product_15(8) <= '0';
partial_product_15(9) <= '0';
partial_product_15(10) <= '0';
partial_product_15(11) <= '0';
partial_product_15(12) <= '0';
partial_product_15(13) <= '0';
partial_product_15(14) <= '0';
partial_product_15(15) <= '0';
partial_product_15(16) <= '0';
partial_product_15(17) <= '0';
partial_product_15(18) <= '0';
partial_product_15(19) <= '0';
partial_product_15(20) <= '0';
partial_product_15(21) <= '0';
partial_product_15(22) <= '0';
partial_product_15(23) <= '0';
partial_product_15(24) <= '0';
partial_product_15(25) <= '0';
partial_product_15(26) <= '0';
partial_product_15(27) <= '0';
partial_product_15(28) <= '0';
partial_product_15(29) <= '0';
partial_product_15(30) <= '0';
partial_product_15(31) <= '0';
partial_product_15(32) <= '0';
partial_product_15(33) <= '0';
partial_product_15(34) <= '0';
partial_product_15(35) <= '0';
partial_product_15(36) <= '0';
partial_product_15(37) <= '0';
partial_product_15(38) <= '0';
partial_product_15(39) <= '0';
partial_product_15(40) <= '0';
partial_product_15(41) <= '0';
partial_product_15(42) <= '0';
partial_product_15(43) <= '0';
partial_product_15(44) <= '0';
partial_product_15(45) <= '0';
partial_product_15(46) <= '0';
partial_product_15(47) <= '0';
partial_product_15(48) <= '0';
partial_product_15(49) <= '0';
partial_product_15(50) <= '0';
partial_product_15(51) <= '0';
partial_product_15(52) <= '0';
partial_product_15(53) <= '0';
partial_product_15(54) <= '0';
partial_product_15(55) <= '0';
partial_product_15(56) <= '0';
partial_product_15(57) <= '0';
partial_product_15(58) <= '0';
partial_product_15(59) <= '0';
partial_product_15(60) <= '0';
partial_product_15(61) <= '0';
partial_product_15(62) <= '0';
partial_product_15(63) <= '0';
partial_product_15(64) <= '0';
partial_product_15(65) <= '0';
partial_product_15(66) <= '0';
partial_product_15(67) <= '0';
partial_product_15(68) <= '0';
partial_product_15(69) <= '0';
partial_product_15(70) <= '0';
partial_product_15(71) <= '0';
partial_product_15(72) <= '0';
partial_product_15(73) <= '0';
partial_product_15(74) <= '0';
partial_product_15(75) <= '0';
partial_product_15(76) <= '0';
partial_product_15(77) <= '0';
partial_product_15(78) <= '0';
partial_product_15(79) <= '0';
partial_product_15(80) <= '0';
partial_product_15(81) <= '0';
partial_product_15(82) <= '0';
partial_product_15(83) <= '0';
partial_product_15(84) <= '0';
partial_product_15(85) <= '0';
partial_product_15(86) <= '0';
partial_product_15(87) <= '0';
partial_product_15(88) <= '0';
partial_product_15(89) <= '0';
partial_product_15(90) <= '0';
partial_product_15(91) <= '0';
partial_product_15(92) <= '0';
partial_product_15(93) <= '0';
partial_product_15(94) <= '0';
partial_product_15(95) <= '0';
partial_product_15(96) <= '0';
partial_product_15(97) <= '0';
partial_product_15(98) <= '0';
partial_product_15(99) <= '0';
partial_product_15(100) <= '0';
partial_product_15(101) <= '0';
partial_product_15(102) <= '0';
partial_product_15(103) <= '0';
partial_product_15(104) <= '0';
partial_product_15(105) <= '0';
partial_product_15(106) <= '0';
partial_product_15(107) <= '0';
partial_product_15(108) <= '0';
partial_product_15(109) <= '0';
partial_product_15(110) <= '0';
partial_product_15(111) <= '0';
partial_product_15(112) <= '0';
partial_product_15(113) <= '0';
partial_product_15(114) <= '0';
partial_product_15(115) <= '0';
partial_product_15(116) <= '0';
partial_product_15(117) <= '0';
partial_product_15(118) <= '0';
partial_product_15(119) <= '0';
partial_product_15(120) <= '0';
partial_product_15(121) <= '0';
partial_product_15(122) <= '0';
partial_product_15(123) <= '0';
partial_product_15(124) <= '0';
partial_product_15(125) <= '0';
partial_product_15(126) <= '0';
partial_product_15(127) <= '0';
partial_product_15(128) <= '0';
partial_product_15(129) <= '0';
partial_product_15(130) <= '0';
partial_product_15(131) <= '0';
partial_product_15(132) <= '0';
partial_product_15(133) <= '0';
partial_product_15(134) <= '0';
partial_product_15(135) <= '0';
partial_product_15(136) <= '0';
partial_product_15(137) <= '0';
partial_product_15(138) <= '0';
partial_product_15(139) <= '0';
partial_product_15(140) <= '0';
partial_product_15(141) <= '0';
partial_product_15(142) <= '0';
partial_product_15(143) <= '0';
partial_product_15(144) <= '0';
partial_product_15(145) <= '0';
partial_product_15(146) <= '0';
partial_product_15(147) <= '0';
partial_product_15(148) <= '0';
partial_product_15(149) <= '0';
partial_product_15(150) <= '0';
partial_product_15(151) <= '0';
partial_product_15(152) <= '0';
partial_product_15(153) <= temp_mult_81(153);
partial_product_15(154) <= temp_mult_81(154);
partial_product_15(155) <= temp_mult_81(155);
partial_product_15(156) <= temp_mult_81(156);
partial_product_15(157) <= temp_mult_81(157);
partial_product_15(158) <= temp_mult_81(158);
partial_product_15(159) <= temp_mult_81(159);
partial_product_15(160) <= temp_mult_81(160);
partial_product_15(161) <= temp_mult_81(161);
partial_product_15(162) <= temp_mult_81(162);
partial_product_15(163) <= temp_mult_81(163);
partial_product_15(164) <= temp_mult_81(164);
partial_product_15(165) <= temp_mult_81(165);
partial_product_15(166) <= temp_mult_81(166);
partial_product_15(167) <= temp_mult_81(167);
partial_product_15(168) <= temp_mult_81(168);
partial_product_15(169) <= temp_mult_81(169);
partial_product_15(170) <= temp_mult_81(170);
partial_product_15(171) <= temp_mult_81(171);
partial_product_15(172) <= temp_mult_81(172);
partial_product_15(173) <= temp_mult_81(173);
partial_product_15(174) <= temp_mult_81(174);
partial_product_15(175) <= temp_mult_81(175);
partial_product_15(176) <= temp_mult_81(176);
partial_product_15(177) <= temp_mult_81(177);
partial_product_15(178) <= temp_mult_81(178);
partial_product_15(179) <= temp_mult_81(179);
partial_product_15(180) <= temp_mult_81(180);
partial_product_15(181) <= temp_mult_81(181);
partial_product_15(182) <= temp_mult_81(182);
partial_product_15(183) <= temp_mult_81(183);
partial_product_15(184) <= temp_mult_81(184);
partial_product_15(185) <= temp_mult_81(185);
partial_product_15(186) <= temp_mult_81(186);
partial_product_15(187) <= temp_mult_81(187);
partial_product_15(188) <= temp_mult_81(188);
partial_product_15(189) <= temp_mult_81(189);
partial_product_15(190) <= temp_mult_81(190);
partial_product_15(191) <= temp_mult_81(191);
partial_product_15(192) <= temp_mult_81(192);
partial_product_15(193) <= temp_mult_81(193);
partial_product_15(194) <= temp_mult_90(194);
partial_product_15(195) <= temp_mult_90(195);
partial_product_15(196) <= temp_mult_90(196);
partial_product_15(197) <= temp_mult_90(197);
partial_product_15(198) <= temp_mult_90(198);
partial_product_15(199) <= temp_mult_90(199);
partial_product_15(200) <= temp_mult_90(200);
partial_product_15(201) <= temp_mult_90(201);
partial_product_15(202) <= temp_mult_90(202);
partial_product_15(203) <= temp_mult_90(203);
partial_product_15(204) <= temp_mult_90(204);
partial_product_15(205) <= temp_mult_90(205);
partial_product_15(206) <= temp_mult_90(206);
partial_product_15(207) <= temp_mult_90(207);
partial_product_15(208) <= temp_mult_90(208);
partial_product_15(209) <= temp_mult_90(209);
partial_product_15(210) <= temp_mult_90(210);
partial_product_15(211) <= temp_mult_90(211);
partial_product_15(212) <= temp_mult_90(212);
partial_product_15(213) <= temp_mult_90(213);
partial_product_15(214) <= temp_mult_90(214);
partial_product_15(215) <= temp_mult_90(215);
partial_product_15(216) <= temp_mult_90(216);
partial_product_15(217) <= temp_mult_90(217);
partial_product_15(218) <= temp_mult_90(218);
partial_product_15(219) <= temp_mult_90(219);
partial_product_15(220) <= temp_mult_90(220);
partial_product_15(221) <= temp_mult_90(221);
partial_product_15(222) <= temp_mult_90(222);
partial_product_15(223) <= temp_mult_90(223);
partial_product_15(224) <= temp_mult_90(224);
partial_product_15(225) <= temp_mult_90(225);
partial_product_15(226) <= temp_mult_90(226);
partial_product_15(227) <= temp_mult_90(227);
partial_product_15(228) <= temp_mult_90(228);
partial_product_15(229) <= temp_mult_90(229);
partial_product_15(230) <= temp_mult_90(230);
partial_product_15(231) <= temp_mult_90(231);
partial_product_15(232) <= temp_mult_90(232);
partial_product_15(233) <= temp_mult_90(233);
partial_product_15(234) <= temp_mult_90(234);
partial_product_15(235) <= temp_mult_99(235);
partial_product_15(236) <= temp_mult_99(236);
partial_product_15(237) <= temp_mult_99(237);
partial_product_15(238) <= temp_mult_99(238);
partial_product_15(239) <= temp_mult_99(239);
partial_product_15(240) <= temp_mult_99(240);
partial_product_15(241) <= temp_mult_99(241);
partial_product_15(242) <= temp_mult_99(242);
partial_product_15(243) <= temp_mult_99(243);
partial_product_15(244) <= temp_mult_99(244);
partial_product_15(245) <= temp_mult_99(245);
partial_product_15(246) <= temp_mult_99(246);
partial_product_15(247) <= temp_mult_99(247);
partial_product_15(248) <= temp_mult_99(248);
partial_product_15(249) <= temp_mult_99(249);
partial_product_15(250) <= temp_mult_99(250);
partial_product_15(251) <= temp_mult_99(251);
partial_product_15(252) <= temp_mult_99(252);
partial_product_15(253) <= temp_mult_99(253);
partial_product_15(254) <= temp_mult_99(254);
partial_product_15(255) <= temp_mult_99(255);
partial_product_15(256) <= temp_mult_99(256);
partial_product_15(257) <= temp_mult_99(257);
partial_product_15(258) <= temp_mult_99(258);
partial_product_15(259) <= temp_mult_99(259);
partial_product_15(260) <= temp_mult_99(260);
partial_product_15(261) <= temp_mult_99(261);
partial_product_15(262) <= temp_mult_99(262);
partial_product_15(263) <= temp_mult_99(263);
partial_product_15(264) <= temp_mult_99(264);
partial_product_15(265) <= temp_mult_99(265);
partial_product_15(266) <= temp_mult_99(266);
partial_product_15(267) <= temp_mult_99(267);
partial_product_15(268) <= temp_mult_99(268);
partial_product_15(269) <= temp_mult_99(269);
partial_product_15(270) <= temp_mult_99(270);
partial_product_15(271) <= temp_mult_99(271);
partial_product_15(272) <= temp_mult_99(272);
partial_product_15(273) <= temp_mult_99(273);
partial_product_15(274) <= temp_mult_99(274);
partial_product_15(275) <= temp_mult_99(275);
partial_product_15(276) <= temp_mult_108(276);
partial_product_15(277) <= temp_mult_108(277);
partial_product_15(278) <= temp_mult_108(278);
partial_product_15(279) <= temp_mult_108(279);
partial_product_15(280) <= temp_mult_108(280);
partial_product_15(281) <= temp_mult_108(281);
partial_product_15(282) <= temp_mult_108(282);
partial_product_15(283) <= temp_mult_108(283);
partial_product_15(284) <= temp_mult_108(284);
partial_product_15(285) <= temp_mult_108(285);
partial_product_15(286) <= temp_mult_108(286);
partial_product_15(287) <= temp_mult_108(287);
partial_product_15(288) <= temp_mult_108(288);
partial_product_15(289) <= temp_mult_108(289);
partial_product_15(290) <= temp_mult_108(290);
partial_product_15(291) <= temp_mult_108(291);
partial_product_15(292) <= temp_mult_108(292);
partial_product_15(293) <= temp_mult_108(293);
partial_product_15(294) <= temp_mult_108(294);
partial_product_15(295) <= temp_mult_108(295);
partial_product_15(296) <= temp_mult_108(296);
partial_product_15(297) <= temp_mult_108(297);
partial_product_15(298) <= temp_mult_108(298);
partial_product_15(299) <= temp_mult_108(299);
partial_product_15(300) <= temp_mult_108(300);
partial_product_15(301) <= temp_mult_108(301);
partial_product_15(302) <= temp_mult_108(302);
partial_product_15(303) <= temp_mult_108(303);
partial_product_15(304) <= temp_mult_108(304);
partial_product_15(305) <= temp_mult_108(305);
partial_product_15(306) <= temp_mult_108(306);
partial_product_15(307) <= temp_mult_108(307);
partial_product_15(308) <= temp_mult_108(308);
partial_product_15(309) <= temp_mult_108(309);
partial_product_15(310) <= temp_mult_108(310);
partial_product_15(311) <= temp_mult_108(311);
partial_product_15(312) <= temp_mult_108(312);
partial_product_15(313) <= temp_mult_108(313);
partial_product_15(314) <= temp_mult_108(314);
partial_product_15(315) <= temp_mult_108(315);
partial_product_15(316) <= temp_mult_108(316);
partial_product_15(317) <= temp_mult_117(317);
partial_product_15(318) <= temp_mult_117(318);
partial_product_15(319) <= temp_mult_117(319);
partial_product_15(320) <= temp_mult_117(320);
partial_product_15(321) <= temp_mult_117(321);
partial_product_15(322) <= temp_mult_117(322);
partial_product_15(323) <= temp_mult_117(323);
partial_product_15(324) <= temp_mult_117(324);
partial_product_15(325) <= temp_mult_117(325);
partial_product_15(326) <= temp_mult_117(326);
partial_product_15(327) <= temp_mult_117(327);
partial_product_15(328) <= temp_mult_117(328);
partial_product_15(329) <= temp_mult_117(329);
partial_product_15(330) <= temp_mult_117(330);
partial_product_15(331) <= temp_mult_117(331);
partial_product_15(332) <= temp_mult_117(332);
partial_product_15(333) <= temp_mult_117(333);
partial_product_15(334) <= temp_mult_117(334);
partial_product_15(335) <= temp_mult_117(335);
partial_product_15(336) <= temp_mult_117(336);
partial_product_15(337) <= temp_mult_117(337);
partial_product_15(338) <= temp_mult_117(338);
partial_product_15(339) <= temp_mult_117(339);
partial_product_15(340) <= temp_mult_117(340);
partial_product_15(341) <= temp_mult_117(341);
partial_product_15(342) <= temp_mult_117(342);
partial_product_15(343) <= temp_mult_117(343);
partial_product_15(344) <= temp_mult_117(344);
partial_product_15(345) <= temp_mult_117(345);
partial_product_15(346) <= temp_mult_117(346);
partial_product_15(347) <= temp_mult_117(347);
partial_product_15(348) <= temp_mult_117(348);
partial_product_15(349) <= temp_mult_117(349);
partial_product_15(350) <= temp_mult_117(350);
partial_product_15(351) <= temp_mult_117(351);
partial_product_15(352) <= temp_mult_117(352);
partial_product_15(353) <= temp_mult_117(353);
partial_product_15(354) <= temp_mult_117(354);
partial_product_15(355) <= temp_mult_117(355);
partial_product_15(356) <= temp_mult_117(356);
partial_product_15(357) <= temp_mult_117(357);
partial_product_15(358) <= '0';
partial_product_15(359) <= '0';
partial_product_15(360) <= '0';
partial_product_15(361) <= '0';
partial_product_15(362) <= '0';
partial_product_15(363) <= '0';
partial_product_15(364) <= '0';
partial_product_15(365) <= '0';
partial_product_15(366) <= '0';
partial_product_15(367) <= '0';
partial_product_15(368) <= '0';
partial_product_15(369) <= '0';
partial_product_15(370) <= '0';
partial_product_15(371) <= '0';
partial_product_15(372) <= '0';
partial_product_15(373) <= '0';
partial_product_15(374) <= '0';
partial_product_15(375) <= '0';
partial_product_15(376) <= '0';
partial_product_15(377) <= '0';
partial_product_15(378) <= '0';
partial_product_15(379) <= '0';
partial_product_15(380) <= '0';
partial_product_15(381) <= '0';
partial_product_15(382) <= '0';
partial_product_15(383) <= '0';
partial_product_15(384) <= '0';
partial_product_15(385) <= '0';
partial_product_15(386) <= '0';
partial_product_15(387) <= '0';
partial_product_15(388) <= '0';
partial_product_15(389) <= '0';
partial_product_15(390) <= '0';
partial_product_15(391) <= '0';
partial_product_15(392) <= '0';
partial_product_15(393) <= '0';
partial_product_15(394) <= '0';
partial_product_15(395) <= '0';
partial_product_15(396) <= '0';
partial_product_15(397) <= '0';
partial_product_15(398) <= '0';
partial_product_15(399) <= '0';
partial_product_15(400) <= '0';
partial_product_15(401) <= '0';
partial_product_15(402) <= '0';
partial_product_15(403) <= '0';
partial_product_15(404) <= '0';
partial_product_15(405) <= '0';
partial_product_15(406) <= '0';
partial_product_15(407) <= '0';
partial_product_15(408) <= '0';
partial_product_15(409) <= '0';
partial_product_15(410) <= '0';
partial_product_15(411) <= '0';
partial_product_15(412) <= '0';
partial_product_15(413) <= '0';
partial_product_15(414) <= '0';
partial_product_15(415) <= '0';
partial_product_15(416) <= '0';
partial_product_15(417) <= '0';
partial_product_15(418) <= '0';
partial_product_15(419) <= '0';
partial_product_15(420) <= '0';
partial_product_15(421) <= '0';
partial_product_15(422) <= '0';
partial_product_15(423) <= '0';
partial_product_15(424) <= '0';
partial_product_15(425) <= '0';
partial_product_15(426) <= '0';
partial_product_15(427) <= '0';
partial_product_15(428) <= '0';
partial_product_15(429) <= '0';
partial_product_15(430) <= '0';
partial_product_15(431) <= '0';
partial_product_15(432) <= '0';
partial_product_15(433) <= '0';
partial_product_15(434) <= '0';
partial_product_15(435) <= '0';
partial_product_15(436) <= '0';
partial_product_15(437) <= '0';
partial_product_15(438) <= '0';
partial_product_15(439) <= '0';
partial_product_15(440) <= '0';
partial_product_15(441) <= '0';
partial_product_15(442) <= '0';
partial_product_15(443) <= '0';
partial_product_15(444) <= '0';
partial_product_15(445) <= '0';
partial_product_15(446) <= '0';
partial_product_15(447) <= '0';
partial_product_15(448) <= '0';
partial_product_15(449) <= '0';
partial_product_15(450) <= '0';
partial_product_15(451) <= '0';
partial_product_15(452) <= '0';
partial_product_15(453) <= '0';
partial_product_15(454) <= '0';
partial_product_15(455) <= '0';
partial_product_15(456) <= '0';
partial_product_15(457) <= '0';
partial_product_15(458) <= '0';
partial_product_15(459) <= '0';
partial_product_15(460) <= '0';
partial_product_15(461) <= '0';
partial_product_15(462) <= '0';
partial_product_15(463) <= '0';
partial_product_15(464) <= '0';
partial_product_15(465) <= '0';
partial_product_15(466) <= '0';
partial_product_15(467) <= '0';
partial_product_15(468) <= '0';
partial_product_15(469) <= '0';
partial_product_15(470) <= '0';
partial_product_15(471) <= '0';
partial_product_15(472) <= '0';
partial_product_15(473) <= '0';
partial_product_15(474) <= '0';
partial_product_15(475) <= '0';
partial_product_15(476) <= '0';
partial_product_15(477) <= '0';
partial_product_15(478) <= '0';
partial_product_15(479) <= '0';
partial_product_15(480) <= '0';
partial_product_15(481) <= '0';
partial_product_15(482) <= '0';
partial_product_15(483) <= '0';
partial_product_15(484) <= '0';
partial_product_15(485) <= '0';
partial_product_15(486) <= '0';
partial_product_15(487) <= '0';
partial_product_15(488) <= '0';
partial_product_15(489) <= '0';
partial_product_15(490) <= '0';
partial_product_15(491) <= '0';
partial_product_15(492) <= '0';
partial_product_15(493) <= '0';
partial_product_15(494) <= '0';
partial_product_15(495) <= '0';
partial_product_15(496) <= '0';
partial_product_15(497) <= '0';
partial_product_15(498) <= '0';
partial_product_15(499) <= '0';
partial_product_15(500) <= '0';
partial_product_15(501) <= '0';
partial_product_15(502) <= '0';
partial_product_15(503) <= '0';
partial_product_15(504) <= '0';
partial_product_15(505) <= '0';
partial_product_15(506) <= '0';
partial_product_15(507) <= '0';
partial_product_15(508) <= '0';
partial_product_15(509) <= '0';
partial_product_15(510) <= '0';
partial_product_15(511) <= '0';
partial_product_15(512) <= '0';
partial_product_16(0) <= '0';
partial_product_16(1) <= '0';
partial_product_16(2) <= '0';
partial_product_16(3) <= '0';
partial_product_16(4) <= '0';
partial_product_16(5) <= '0';
partial_product_16(6) <= '0';
partial_product_16(7) <= '0';
partial_product_16(8) <= '0';
partial_product_16(9) <= '0';
partial_product_16(10) <= '0';
partial_product_16(11) <= '0';
partial_product_16(12) <= '0';
partial_product_16(13) <= '0';
partial_product_16(14) <= '0';
partial_product_16(15) <= '0';
partial_product_16(16) <= '0';
partial_product_16(17) <= '0';
partial_product_16(18) <= '0';
partial_product_16(19) <= '0';
partial_product_16(20) <= '0';
partial_product_16(21) <= '0';
partial_product_16(22) <= '0';
partial_product_16(23) <= '0';
partial_product_16(24) <= '0';
partial_product_16(25) <= '0';
partial_product_16(26) <= '0';
partial_product_16(27) <= '0';
partial_product_16(28) <= '0';
partial_product_16(29) <= '0';
partial_product_16(30) <= '0';
partial_product_16(31) <= '0';
partial_product_16(32) <= '0';
partial_product_16(33) <= '0';
partial_product_16(34) <= '0';
partial_product_16(35) <= '0';
partial_product_16(36) <= '0';
partial_product_16(37) <= '0';
partial_product_16(38) <= '0';
partial_product_16(39) <= '0';
partial_product_16(40) <= '0';
partial_product_16(41) <= '0';
partial_product_16(42) <= '0';
partial_product_16(43) <= '0';
partial_product_16(44) <= '0';
partial_product_16(45) <= '0';
partial_product_16(46) <= '0';
partial_product_16(47) <= '0';
partial_product_16(48) <= '0';
partial_product_16(49) <= '0';
partial_product_16(50) <= '0';
partial_product_16(51) <= '0';
partial_product_16(52) <= '0';
partial_product_16(53) <= '0';
partial_product_16(54) <= '0';
partial_product_16(55) <= '0';
partial_product_16(56) <= '0';
partial_product_16(57) <= '0';
partial_product_16(58) <= '0';
partial_product_16(59) <= '0';
partial_product_16(60) <= '0';
partial_product_16(61) <= '0';
partial_product_16(62) <= '0';
partial_product_16(63) <= '0';
partial_product_16(64) <= '0';
partial_product_16(65) <= '0';
partial_product_16(66) <= '0';
partial_product_16(67) <= '0';
partial_product_16(68) <= '0';
partial_product_16(69) <= '0';
partial_product_16(70) <= '0';
partial_product_16(71) <= '0';
partial_product_16(72) <= '0';
partial_product_16(73) <= '0';
partial_product_16(74) <= '0';
partial_product_16(75) <= '0';
partial_product_16(76) <= '0';
partial_product_16(77) <= '0';
partial_product_16(78) <= '0';
partial_product_16(79) <= '0';
partial_product_16(80) <= '0';
partial_product_16(81) <= '0';
partial_product_16(82) <= '0';
partial_product_16(83) <= '0';
partial_product_16(84) <= '0';
partial_product_16(85) <= '0';
partial_product_16(86) <= '0';
partial_product_16(87) <= '0';
partial_product_16(88) <= '0';
partial_product_16(89) <= '0';
partial_product_16(90) <= '0';
partial_product_16(91) <= '0';
partial_product_16(92) <= '0';
partial_product_16(93) <= '0';
partial_product_16(94) <= '0';
partial_product_16(95) <= '0';
partial_product_16(96) <= '0';
partial_product_16(97) <= '0';
partial_product_16(98) <= '0';
partial_product_16(99) <= '0';
partial_product_16(100) <= '0';
partial_product_16(101) <= '0';
partial_product_16(102) <= '0';
partial_product_16(103) <= '0';
partial_product_16(104) <= '0';
partial_product_16(105) <= '0';
partial_product_16(106) <= '0';
partial_product_16(107) <= '0';
partial_product_16(108) <= '0';
partial_product_16(109) <= '0';
partial_product_16(110) <= '0';
partial_product_16(111) <= '0';
partial_product_16(112) <= '0';
partial_product_16(113) <= '0';
partial_product_16(114) <= '0';
partial_product_16(115) <= '0';
partial_product_16(116) <= '0';
partial_product_16(117) <= '0';
partial_product_16(118) <= '0';
partial_product_16(119) <= '0';
partial_product_16(120) <= '0';
partial_product_16(121) <= '0';
partial_product_16(122) <= '0';
partial_product_16(123) <= '0';
partial_product_16(124) <= '0';
partial_product_16(125) <= '0';
partial_product_16(126) <= '0';
partial_product_16(127) <= '0';
partial_product_16(128) <= '0';
partial_product_16(129) <= '0';
partial_product_16(130) <= '0';
partial_product_16(131) <= '0';
partial_product_16(132) <= '0';
partial_product_16(133) <= '0';
partial_product_16(134) <= '0';
partial_product_16(135) <= '0';
partial_product_16(136) <= '0';
partial_product_16(137) <= '0';
partial_product_16(138) <= '0';
partial_product_16(139) <= '0';
partial_product_16(140) <= '0';
partial_product_16(141) <= '0';
partial_product_16(142) <= '0';
partial_product_16(143) <= '0';
partial_product_16(144) <= '0';
partial_product_16(145) <= '0';
partial_product_16(146) <= '0';
partial_product_16(147) <= '0';
partial_product_16(148) <= '0';
partial_product_16(149) <= '0';
partial_product_16(150) <= '0';
partial_product_16(151) <= '0';
partial_product_16(152) <= '0';
partial_product_16(153) <= '0';
partial_product_16(154) <= '0';
partial_product_16(155) <= '0';
partial_product_16(156) <= '0';
partial_product_16(157) <= '0';
partial_product_16(158) <= '0';
partial_product_16(159) <= '0';
partial_product_16(160) <= '0';
partial_product_16(161) <= '0';
partial_product_16(162) <= '0';
partial_product_16(163) <= '0';
partial_product_16(164) <= '0';
partial_product_16(165) <= '0';
partial_product_16(166) <= '0';
partial_product_16(167) <= '0';
partial_product_16(168) <= temp_mult_56(168);
partial_product_16(169) <= temp_mult_56(169);
partial_product_16(170) <= temp_mult_56(170);
partial_product_16(171) <= temp_mult_56(171);
partial_product_16(172) <= temp_mult_56(172);
partial_product_16(173) <= temp_mult_56(173);
partial_product_16(174) <= temp_mult_56(174);
partial_product_16(175) <= temp_mult_56(175);
partial_product_16(176) <= temp_mult_56(176);
partial_product_16(177) <= temp_mult_56(177);
partial_product_16(178) <= temp_mult_56(178);
partial_product_16(179) <= temp_mult_56(179);
partial_product_16(180) <= temp_mult_56(180);
partial_product_16(181) <= temp_mult_56(181);
partial_product_16(182) <= temp_mult_56(182);
partial_product_16(183) <= temp_mult_56(183);
partial_product_16(184) <= temp_mult_56(184);
partial_product_16(185) <= temp_mult_56(185);
partial_product_16(186) <= temp_mult_56(186);
partial_product_16(187) <= temp_mult_56(187);
partial_product_16(188) <= temp_mult_56(188);
partial_product_16(189) <= temp_mult_56(189);
partial_product_16(190) <= temp_mult_56(190);
partial_product_16(191) <= temp_mult_56(191);
partial_product_16(192) <= temp_mult_56(192);
partial_product_16(193) <= temp_mult_56(193);
partial_product_16(194) <= temp_mult_56(194);
partial_product_16(195) <= temp_mult_56(195);
partial_product_16(196) <= temp_mult_56(196);
partial_product_16(197) <= temp_mult_56(197);
partial_product_16(198) <= temp_mult_56(198);
partial_product_16(199) <= temp_mult_56(199);
partial_product_16(200) <= temp_mult_56(200);
partial_product_16(201) <= temp_mult_56(201);
partial_product_16(202) <= temp_mult_56(202);
partial_product_16(203) <= temp_mult_56(203);
partial_product_16(204) <= temp_mult_56(204);
partial_product_16(205) <= temp_mult_56(205);
partial_product_16(206) <= temp_mult_56(206);
partial_product_16(207) <= temp_mult_56(207);
partial_product_16(208) <= temp_mult_56(208);
partial_product_16(209) <= temp_mult_65(209);
partial_product_16(210) <= temp_mult_65(210);
partial_product_16(211) <= temp_mult_65(211);
partial_product_16(212) <= temp_mult_65(212);
partial_product_16(213) <= temp_mult_65(213);
partial_product_16(214) <= temp_mult_65(214);
partial_product_16(215) <= temp_mult_65(215);
partial_product_16(216) <= temp_mult_65(216);
partial_product_16(217) <= temp_mult_65(217);
partial_product_16(218) <= temp_mult_65(218);
partial_product_16(219) <= temp_mult_65(219);
partial_product_16(220) <= temp_mult_65(220);
partial_product_16(221) <= temp_mult_65(221);
partial_product_16(222) <= temp_mult_65(222);
partial_product_16(223) <= temp_mult_65(223);
partial_product_16(224) <= temp_mult_65(224);
partial_product_16(225) <= temp_mult_65(225);
partial_product_16(226) <= temp_mult_65(226);
partial_product_16(227) <= temp_mult_65(227);
partial_product_16(228) <= temp_mult_65(228);
partial_product_16(229) <= temp_mult_65(229);
partial_product_16(230) <= temp_mult_65(230);
partial_product_16(231) <= temp_mult_65(231);
partial_product_16(232) <= temp_mult_65(232);
partial_product_16(233) <= temp_mult_65(233);
partial_product_16(234) <= temp_mult_65(234);
partial_product_16(235) <= temp_mult_65(235);
partial_product_16(236) <= temp_mult_65(236);
partial_product_16(237) <= temp_mult_65(237);
partial_product_16(238) <= temp_mult_65(238);
partial_product_16(239) <= temp_mult_65(239);
partial_product_16(240) <= temp_mult_65(240);
partial_product_16(241) <= temp_mult_65(241);
partial_product_16(242) <= temp_mult_65(242);
partial_product_16(243) <= temp_mult_65(243);
partial_product_16(244) <= temp_mult_65(244);
partial_product_16(245) <= temp_mult_65(245);
partial_product_16(246) <= temp_mult_65(246);
partial_product_16(247) <= temp_mult_65(247);
partial_product_16(248) <= temp_mult_65(248);
partial_product_16(249) <= temp_mult_65(249);
partial_product_16(250) <= temp_mult_74(250);
partial_product_16(251) <= temp_mult_74(251);
partial_product_16(252) <= temp_mult_74(252);
partial_product_16(253) <= temp_mult_74(253);
partial_product_16(254) <= temp_mult_74(254);
partial_product_16(255) <= temp_mult_74(255);
partial_product_16(256) <= temp_mult_74(256);
partial_product_16(257) <= temp_mult_74(257);
partial_product_16(258) <= temp_mult_74(258);
partial_product_16(259) <= temp_mult_74(259);
partial_product_16(260) <= temp_mult_74(260);
partial_product_16(261) <= temp_mult_74(261);
partial_product_16(262) <= temp_mult_74(262);
partial_product_16(263) <= temp_mult_74(263);
partial_product_16(264) <= temp_mult_74(264);
partial_product_16(265) <= temp_mult_74(265);
partial_product_16(266) <= temp_mult_74(266);
partial_product_16(267) <= temp_mult_74(267);
partial_product_16(268) <= temp_mult_74(268);
partial_product_16(269) <= temp_mult_74(269);
partial_product_16(270) <= temp_mult_74(270);
partial_product_16(271) <= temp_mult_74(271);
partial_product_16(272) <= temp_mult_74(272);
partial_product_16(273) <= temp_mult_74(273);
partial_product_16(274) <= temp_mult_74(274);
partial_product_16(275) <= temp_mult_74(275);
partial_product_16(276) <= temp_mult_74(276);
partial_product_16(277) <= temp_mult_74(277);
partial_product_16(278) <= temp_mult_74(278);
partial_product_16(279) <= temp_mult_74(279);
partial_product_16(280) <= temp_mult_74(280);
partial_product_16(281) <= temp_mult_74(281);
partial_product_16(282) <= temp_mult_74(282);
partial_product_16(283) <= temp_mult_74(283);
partial_product_16(284) <= temp_mult_74(284);
partial_product_16(285) <= temp_mult_74(285);
partial_product_16(286) <= temp_mult_74(286);
partial_product_16(287) <= temp_mult_74(287);
partial_product_16(288) <= temp_mult_74(288);
partial_product_16(289) <= temp_mult_74(289);
partial_product_16(290) <= temp_mult_74(290);
partial_product_16(291) <= '0';
partial_product_16(292) <= '0';
partial_product_16(293) <= temp_mult_109(293);
partial_product_16(294) <= temp_mult_109(294);
partial_product_16(295) <= temp_mult_109(295);
partial_product_16(296) <= temp_mult_109(296);
partial_product_16(297) <= temp_mult_109(297);
partial_product_16(298) <= temp_mult_109(298);
partial_product_16(299) <= temp_mult_109(299);
partial_product_16(300) <= temp_mult_109(300);
partial_product_16(301) <= temp_mult_109(301);
partial_product_16(302) <= temp_mult_109(302);
partial_product_16(303) <= temp_mult_109(303);
partial_product_16(304) <= temp_mult_109(304);
partial_product_16(305) <= temp_mult_109(305);
partial_product_16(306) <= temp_mult_109(306);
partial_product_16(307) <= temp_mult_109(307);
partial_product_16(308) <= temp_mult_109(308);
partial_product_16(309) <= temp_mult_109(309);
partial_product_16(310) <= temp_mult_109(310);
partial_product_16(311) <= temp_mult_109(311);
partial_product_16(312) <= temp_mult_109(312);
partial_product_16(313) <= temp_mult_109(313);
partial_product_16(314) <= temp_mult_109(314);
partial_product_16(315) <= temp_mult_109(315);
partial_product_16(316) <= temp_mult_109(316);
partial_product_16(317) <= temp_mult_109(317);
partial_product_16(318) <= temp_mult_109(318);
partial_product_16(319) <= temp_mult_109(319);
partial_product_16(320) <= temp_mult_109(320);
partial_product_16(321) <= temp_mult_109(321);
partial_product_16(322) <= temp_mult_109(322);
partial_product_16(323) <= temp_mult_109(323);
partial_product_16(324) <= temp_mult_109(324);
partial_product_16(325) <= temp_mult_109(325);
partial_product_16(326) <= temp_mult_109(326);
partial_product_16(327) <= temp_mult_109(327);
partial_product_16(328) <= temp_mult_109(328);
partial_product_16(329) <= temp_mult_109(329);
partial_product_16(330) <= temp_mult_109(330);
partial_product_16(331) <= temp_mult_109(331);
partial_product_16(332) <= temp_mult_109(332);
partial_product_16(333) <= temp_mult_109(333);
partial_product_16(334) <= temp_mult_118(334);
partial_product_16(335) <= temp_mult_118(335);
partial_product_16(336) <= temp_mult_118(336);
partial_product_16(337) <= temp_mult_118(337);
partial_product_16(338) <= temp_mult_118(338);
partial_product_16(339) <= temp_mult_118(339);
partial_product_16(340) <= temp_mult_118(340);
partial_product_16(341) <= temp_mult_118(341);
partial_product_16(342) <= temp_mult_118(342);
partial_product_16(343) <= temp_mult_118(343);
partial_product_16(344) <= temp_mult_118(344);
partial_product_16(345) <= temp_mult_118(345);
partial_product_16(346) <= temp_mult_118(346);
partial_product_16(347) <= temp_mult_118(347);
partial_product_16(348) <= temp_mult_118(348);
partial_product_16(349) <= temp_mult_118(349);
partial_product_16(350) <= temp_mult_118(350);
partial_product_16(351) <= temp_mult_118(351);
partial_product_16(352) <= temp_mult_118(352);
partial_product_16(353) <= temp_mult_118(353);
partial_product_16(354) <= temp_mult_118(354);
partial_product_16(355) <= temp_mult_118(355);
partial_product_16(356) <= temp_mult_118(356);
partial_product_16(357) <= temp_mult_118(357);
partial_product_16(358) <= temp_mult_118(358);
partial_product_16(359) <= temp_mult_118(359);
partial_product_16(360) <= temp_mult_118(360);
partial_product_16(361) <= temp_mult_118(361);
partial_product_16(362) <= temp_mult_118(362);
partial_product_16(363) <= temp_mult_118(363);
partial_product_16(364) <= temp_mult_118(364);
partial_product_16(365) <= temp_mult_118(365);
partial_product_16(366) <= temp_mult_118(366);
partial_product_16(367) <= temp_mult_118(367);
partial_product_16(368) <= temp_mult_118(368);
partial_product_16(369) <= temp_mult_118(369);
partial_product_16(370) <= temp_mult_118(370);
partial_product_16(371) <= temp_mult_118(371);
partial_product_16(372) <= temp_mult_118(372);
partial_product_16(373) <= temp_mult_118(373);
partial_product_16(374) <= temp_mult_118(374);
partial_product_16(375) <= '0';
partial_product_16(376) <= '0';
partial_product_16(377) <= '0';
partial_product_16(378) <= '0';
partial_product_16(379) <= '0';
partial_product_16(380) <= '0';
partial_product_16(381) <= '0';
partial_product_16(382) <= '0';
partial_product_16(383) <= '0';
partial_product_16(384) <= '0';
partial_product_16(385) <= '0';
partial_product_16(386) <= '0';
partial_product_16(387) <= '0';
partial_product_16(388) <= '0';
partial_product_16(389) <= '0';
partial_product_16(390) <= '0';
partial_product_16(391) <= '0';
partial_product_16(392) <= '0';
partial_product_16(393) <= '0';
partial_product_16(394) <= '0';
partial_product_16(395) <= '0';
partial_product_16(396) <= '0';
partial_product_16(397) <= '0';
partial_product_16(398) <= '0';
partial_product_16(399) <= '0';
partial_product_16(400) <= '0';
partial_product_16(401) <= '0';
partial_product_16(402) <= '0';
partial_product_16(403) <= '0';
partial_product_16(404) <= '0';
partial_product_16(405) <= '0';
partial_product_16(406) <= '0';
partial_product_16(407) <= '0';
partial_product_16(408) <= '0';
partial_product_16(409) <= '0';
partial_product_16(410) <= '0';
partial_product_16(411) <= '0';
partial_product_16(412) <= '0';
partial_product_16(413) <= '0';
partial_product_16(414) <= '0';
partial_product_16(415) <= '0';
partial_product_16(416) <= '0';
partial_product_16(417) <= '0';
partial_product_16(418) <= '0';
partial_product_16(419) <= '0';
partial_product_16(420) <= '0';
partial_product_16(421) <= '0';
partial_product_16(422) <= '0';
partial_product_16(423) <= '0';
partial_product_16(424) <= '0';
partial_product_16(425) <= '0';
partial_product_16(426) <= '0';
partial_product_16(427) <= '0';
partial_product_16(428) <= '0';
partial_product_16(429) <= '0';
partial_product_16(430) <= '0';
partial_product_16(431) <= '0';
partial_product_16(432) <= '0';
partial_product_16(433) <= '0';
partial_product_16(434) <= '0';
partial_product_16(435) <= '0';
partial_product_16(436) <= '0';
partial_product_16(437) <= '0';
partial_product_16(438) <= '0';
partial_product_16(439) <= '0';
partial_product_16(440) <= '0';
partial_product_16(441) <= '0';
partial_product_16(442) <= '0';
partial_product_16(443) <= '0';
partial_product_16(444) <= '0';
partial_product_16(445) <= '0';
partial_product_16(446) <= '0';
partial_product_16(447) <= '0';
partial_product_16(448) <= '0';
partial_product_16(449) <= '0';
partial_product_16(450) <= '0';
partial_product_16(451) <= '0';
partial_product_16(452) <= '0';
partial_product_16(453) <= '0';
partial_product_16(454) <= '0';
partial_product_16(455) <= '0';
partial_product_16(456) <= '0';
partial_product_16(457) <= '0';
partial_product_16(458) <= '0';
partial_product_16(459) <= '0';
partial_product_16(460) <= '0';
partial_product_16(461) <= '0';
partial_product_16(462) <= '0';
partial_product_16(463) <= '0';
partial_product_16(464) <= '0';
partial_product_16(465) <= '0';
partial_product_16(466) <= '0';
partial_product_16(467) <= '0';
partial_product_16(468) <= '0';
partial_product_16(469) <= '0';
partial_product_16(470) <= '0';
partial_product_16(471) <= '0';
partial_product_16(472) <= '0';
partial_product_16(473) <= '0';
partial_product_16(474) <= '0';
partial_product_16(475) <= '0';
partial_product_16(476) <= '0';
partial_product_16(477) <= '0';
partial_product_16(478) <= '0';
partial_product_16(479) <= '0';
partial_product_16(480) <= '0';
partial_product_16(481) <= '0';
partial_product_16(482) <= '0';
partial_product_16(483) <= '0';
partial_product_16(484) <= '0';
partial_product_16(485) <= '0';
partial_product_16(486) <= '0';
partial_product_16(487) <= '0';
partial_product_16(488) <= '0';
partial_product_16(489) <= '0';
partial_product_16(490) <= '0';
partial_product_16(491) <= '0';
partial_product_16(492) <= '0';
partial_product_16(493) <= '0';
partial_product_16(494) <= '0';
partial_product_16(495) <= '0';
partial_product_16(496) <= '0';
partial_product_16(497) <= '0';
partial_product_16(498) <= '0';
partial_product_16(499) <= '0';
partial_product_16(500) <= '0';
partial_product_16(501) <= '0';
partial_product_16(502) <= '0';
partial_product_16(503) <= '0';
partial_product_16(504) <= '0';
partial_product_16(505) <= '0';
partial_product_16(506) <= '0';
partial_product_16(507) <= '0';
partial_product_16(508) <= '0';
partial_product_16(509) <= '0';
partial_product_16(510) <= '0';
partial_product_16(511) <= '0';
partial_product_16(512) <= '0';
partial_product_17(0) <= '0';
partial_product_17(1) <= '0';
partial_product_17(2) <= '0';
partial_product_17(3) <= '0';
partial_product_17(4) <= '0';
partial_product_17(5) <= '0';
partial_product_17(6) <= '0';
partial_product_17(7) <= '0';
partial_product_17(8) <= '0';
partial_product_17(9) <= '0';
partial_product_17(10) <= '0';
partial_product_17(11) <= '0';
partial_product_17(12) <= '0';
partial_product_17(13) <= '0';
partial_product_17(14) <= '0';
partial_product_17(15) <= '0';
partial_product_17(16) <= '0';
partial_product_17(17) <= '0';
partial_product_17(18) <= '0';
partial_product_17(19) <= '0';
partial_product_17(20) <= '0';
partial_product_17(21) <= '0';
partial_product_17(22) <= '0';
partial_product_17(23) <= '0';
partial_product_17(24) <= '0';
partial_product_17(25) <= '0';
partial_product_17(26) <= '0';
partial_product_17(27) <= '0';
partial_product_17(28) <= '0';
partial_product_17(29) <= '0';
partial_product_17(30) <= '0';
partial_product_17(31) <= '0';
partial_product_17(32) <= '0';
partial_product_17(33) <= '0';
partial_product_17(34) <= '0';
partial_product_17(35) <= '0';
partial_product_17(36) <= '0';
partial_product_17(37) <= '0';
partial_product_17(38) <= '0';
partial_product_17(39) <= '0';
partial_product_17(40) <= '0';
partial_product_17(41) <= '0';
partial_product_17(42) <= '0';
partial_product_17(43) <= '0';
partial_product_17(44) <= '0';
partial_product_17(45) <= '0';
partial_product_17(46) <= '0';
partial_product_17(47) <= '0';
partial_product_17(48) <= '0';
partial_product_17(49) <= '0';
partial_product_17(50) <= '0';
partial_product_17(51) <= '0';
partial_product_17(52) <= '0';
partial_product_17(53) <= '0';
partial_product_17(54) <= '0';
partial_product_17(55) <= '0';
partial_product_17(56) <= '0';
partial_product_17(57) <= '0';
partial_product_17(58) <= '0';
partial_product_17(59) <= '0';
partial_product_17(60) <= '0';
partial_product_17(61) <= '0';
partial_product_17(62) <= '0';
partial_product_17(63) <= '0';
partial_product_17(64) <= '0';
partial_product_17(65) <= '0';
partial_product_17(66) <= '0';
partial_product_17(67) <= '0';
partial_product_17(68) <= '0';
partial_product_17(69) <= '0';
partial_product_17(70) <= '0';
partial_product_17(71) <= '0';
partial_product_17(72) <= '0';
partial_product_17(73) <= '0';
partial_product_17(74) <= '0';
partial_product_17(75) <= '0';
partial_product_17(76) <= '0';
partial_product_17(77) <= '0';
partial_product_17(78) <= '0';
partial_product_17(79) <= '0';
partial_product_17(80) <= '0';
partial_product_17(81) <= '0';
partial_product_17(82) <= '0';
partial_product_17(83) <= '0';
partial_product_17(84) <= '0';
partial_product_17(85) <= '0';
partial_product_17(86) <= '0';
partial_product_17(87) <= '0';
partial_product_17(88) <= '0';
partial_product_17(89) <= '0';
partial_product_17(90) <= '0';
partial_product_17(91) <= '0';
partial_product_17(92) <= '0';
partial_product_17(93) <= '0';
partial_product_17(94) <= '0';
partial_product_17(95) <= '0';
partial_product_17(96) <= '0';
partial_product_17(97) <= '0';
partial_product_17(98) <= '0';
partial_product_17(99) <= '0';
partial_product_17(100) <= '0';
partial_product_17(101) <= '0';
partial_product_17(102) <= '0';
partial_product_17(103) <= '0';
partial_product_17(104) <= '0';
partial_product_17(105) <= '0';
partial_product_17(106) <= '0';
partial_product_17(107) <= '0';
partial_product_17(108) <= '0';
partial_product_17(109) <= '0';
partial_product_17(110) <= '0';
partial_product_17(111) <= '0';
partial_product_17(112) <= '0';
partial_product_17(113) <= '0';
partial_product_17(114) <= '0';
partial_product_17(115) <= '0';
partial_product_17(116) <= '0';
partial_product_17(117) <= '0';
partial_product_17(118) <= '0';
partial_product_17(119) <= '0';
partial_product_17(120) <= '0';
partial_product_17(121) <= '0';
partial_product_17(122) <= '0';
partial_product_17(123) <= '0';
partial_product_17(124) <= '0';
partial_product_17(125) <= '0';
partial_product_17(126) <= '0';
partial_product_17(127) <= '0';
partial_product_17(128) <= '0';
partial_product_17(129) <= '0';
partial_product_17(130) <= '0';
partial_product_17(131) <= '0';
partial_product_17(132) <= '0';
partial_product_17(133) <= '0';
partial_product_17(134) <= '0';
partial_product_17(135) <= '0';
partial_product_17(136) <= '0';
partial_product_17(137) <= '0';
partial_product_17(138) <= '0';
partial_product_17(139) <= '0';
partial_product_17(140) <= '0';
partial_product_17(141) <= '0';
partial_product_17(142) <= '0';
partial_product_17(143) <= '0';
partial_product_17(144) <= '0';
partial_product_17(145) <= '0';
partial_product_17(146) <= '0';
partial_product_17(147) <= '0';
partial_product_17(148) <= '0';
partial_product_17(149) <= '0';
partial_product_17(150) <= '0';
partial_product_17(151) <= '0';
partial_product_17(152) <= '0';
partial_product_17(153) <= '0';
partial_product_17(154) <= '0';
partial_product_17(155) <= '0';
partial_product_17(156) <= '0';
partial_product_17(157) <= '0';
partial_product_17(158) <= '0';
partial_product_17(159) <= '0';
partial_product_17(160) <= '0';
partial_product_17(161) <= '0';
partial_product_17(162) <= '0';
partial_product_17(163) <= '0';
partial_product_17(164) <= '0';
partial_product_17(165) <= '0';
partial_product_17(166) <= '0';
partial_product_17(167) <= '0';
partial_product_17(168) <= '0';
partial_product_17(169) <= '0';
partial_product_17(170) <= temp_mult_82(170);
partial_product_17(171) <= temp_mult_82(171);
partial_product_17(172) <= temp_mult_82(172);
partial_product_17(173) <= temp_mult_82(173);
partial_product_17(174) <= temp_mult_82(174);
partial_product_17(175) <= temp_mult_82(175);
partial_product_17(176) <= temp_mult_82(176);
partial_product_17(177) <= temp_mult_82(177);
partial_product_17(178) <= temp_mult_82(178);
partial_product_17(179) <= temp_mult_82(179);
partial_product_17(180) <= temp_mult_82(180);
partial_product_17(181) <= temp_mult_82(181);
partial_product_17(182) <= temp_mult_82(182);
partial_product_17(183) <= temp_mult_82(183);
partial_product_17(184) <= temp_mult_82(184);
partial_product_17(185) <= temp_mult_82(185);
partial_product_17(186) <= temp_mult_82(186);
partial_product_17(187) <= temp_mult_82(187);
partial_product_17(188) <= temp_mult_82(188);
partial_product_17(189) <= temp_mult_82(189);
partial_product_17(190) <= temp_mult_82(190);
partial_product_17(191) <= temp_mult_82(191);
partial_product_17(192) <= temp_mult_82(192);
partial_product_17(193) <= temp_mult_82(193);
partial_product_17(194) <= temp_mult_82(194);
partial_product_17(195) <= temp_mult_82(195);
partial_product_17(196) <= temp_mult_82(196);
partial_product_17(197) <= temp_mult_82(197);
partial_product_17(198) <= temp_mult_82(198);
partial_product_17(199) <= temp_mult_82(199);
partial_product_17(200) <= temp_mult_82(200);
partial_product_17(201) <= temp_mult_82(201);
partial_product_17(202) <= temp_mult_82(202);
partial_product_17(203) <= temp_mult_82(203);
partial_product_17(204) <= temp_mult_82(204);
partial_product_17(205) <= temp_mult_82(205);
partial_product_17(206) <= temp_mult_82(206);
partial_product_17(207) <= temp_mult_82(207);
partial_product_17(208) <= temp_mult_82(208);
partial_product_17(209) <= temp_mult_82(209);
partial_product_17(210) <= temp_mult_82(210);
partial_product_17(211) <= temp_mult_91(211);
partial_product_17(212) <= temp_mult_91(212);
partial_product_17(213) <= temp_mult_91(213);
partial_product_17(214) <= temp_mult_91(214);
partial_product_17(215) <= temp_mult_91(215);
partial_product_17(216) <= temp_mult_91(216);
partial_product_17(217) <= temp_mult_91(217);
partial_product_17(218) <= temp_mult_91(218);
partial_product_17(219) <= temp_mult_91(219);
partial_product_17(220) <= temp_mult_91(220);
partial_product_17(221) <= temp_mult_91(221);
partial_product_17(222) <= temp_mult_91(222);
partial_product_17(223) <= temp_mult_91(223);
partial_product_17(224) <= temp_mult_91(224);
partial_product_17(225) <= temp_mult_91(225);
partial_product_17(226) <= temp_mult_91(226);
partial_product_17(227) <= temp_mult_91(227);
partial_product_17(228) <= temp_mult_91(228);
partial_product_17(229) <= temp_mult_91(229);
partial_product_17(230) <= temp_mult_91(230);
partial_product_17(231) <= temp_mult_91(231);
partial_product_17(232) <= temp_mult_91(232);
partial_product_17(233) <= temp_mult_91(233);
partial_product_17(234) <= temp_mult_91(234);
partial_product_17(235) <= temp_mult_91(235);
partial_product_17(236) <= temp_mult_91(236);
partial_product_17(237) <= temp_mult_91(237);
partial_product_17(238) <= temp_mult_91(238);
partial_product_17(239) <= temp_mult_91(239);
partial_product_17(240) <= temp_mult_91(240);
partial_product_17(241) <= temp_mult_91(241);
partial_product_17(242) <= temp_mult_91(242);
partial_product_17(243) <= temp_mult_91(243);
partial_product_17(244) <= temp_mult_91(244);
partial_product_17(245) <= temp_mult_91(245);
partial_product_17(246) <= temp_mult_91(246);
partial_product_17(247) <= temp_mult_91(247);
partial_product_17(248) <= temp_mult_91(248);
partial_product_17(249) <= temp_mult_91(249);
partial_product_17(250) <= temp_mult_91(250);
partial_product_17(251) <= temp_mult_91(251);
partial_product_17(252) <= temp_mult_100(252);
partial_product_17(253) <= temp_mult_100(253);
partial_product_17(254) <= temp_mult_100(254);
partial_product_17(255) <= temp_mult_100(255);
partial_product_17(256) <= temp_mult_100(256);
partial_product_17(257) <= temp_mult_100(257);
partial_product_17(258) <= temp_mult_100(258);
partial_product_17(259) <= temp_mult_100(259);
partial_product_17(260) <= temp_mult_100(260);
partial_product_17(261) <= temp_mult_100(261);
partial_product_17(262) <= temp_mult_100(262);
partial_product_17(263) <= temp_mult_100(263);
partial_product_17(264) <= temp_mult_100(264);
partial_product_17(265) <= temp_mult_100(265);
partial_product_17(266) <= temp_mult_100(266);
partial_product_17(267) <= temp_mult_100(267);
partial_product_17(268) <= temp_mult_100(268);
partial_product_17(269) <= temp_mult_100(269);
partial_product_17(270) <= temp_mult_100(270);
partial_product_17(271) <= temp_mult_100(271);
partial_product_17(272) <= temp_mult_100(272);
partial_product_17(273) <= temp_mult_100(273);
partial_product_17(274) <= temp_mult_100(274);
partial_product_17(275) <= temp_mult_100(275);
partial_product_17(276) <= temp_mult_100(276);
partial_product_17(277) <= temp_mult_100(277);
partial_product_17(278) <= temp_mult_100(278);
partial_product_17(279) <= temp_mult_100(279);
partial_product_17(280) <= temp_mult_100(280);
partial_product_17(281) <= temp_mult_100(281);
partial_product_17(282) <= temp_mult_100(282);
partial_product_17(283) <= temp_mult_100(283);
partial_product_17(284) <= temp_mult_100(284);
partial_product_17(285) <= temp_mult_100(285);
partial_product_17(286) <= temp_mult_100(286);
partial_product_17(287) <= temp_mult_100(287);
partial_product_17(288) <= temp_mult_100(288);
partial_product_17(289) <= temp_mult_100(289);
partial_product_17(290) <= temp_mult_100(290);
partial_product_17(291) <= temp_mult_100(291);
partial_product_17(292) <= temp_mult_100(292);
partial_product_17(293) <= '0';
partial_product_17(294) <= '0';
partial_product_17(295) <= '0';
partial_product_17(296) <= '0';
partial_product_17(297) <= '0';
partial_product_17(298) <= '0';
partial_product_17(299) <= '0';
partial_product_17(300) <= '0';
partial_product_17(301) <= '0';
partial_product_17(302) <= '0';
partial_product_17(303) <= temp_mult_103(303);
partial_product_17(304) <= temp_mult_103(304);
partial_product_17(305) <= temp_mult_103(305);
partial_product_17(306) <= temp_mult_103(306);
partial_product_17(307) <= temp_mult_103(307);
partial_product_17(308) <= temp_mult_103(308);
partial_product_17(309) <= temp_mult_103(309);
partial_product_17(310) <= temp_mult_103(310);
partial_product_17(311) <= temp_mult_103(311);
partial_product_17(312) <= temp_mult_103(312);
partial_product_17(313) <= temp_mult_103(313);
partial_product_17(314) <= temp_mult_103(314);
partial_product_17(315) <= temp_mult_103(315);
partial_product_17(316) <= temp_mult_103(316);
partial_product_17(317) <= temp_mult_103(317);
partial_product_17(318) <= temp_mult_103(318);
partial_product_17(319) <= temp_mult_103(319);
partial_product_17(320) <= temp_mult_103(320);
partial_product_17(321) <= temp_mult_103(321);
partial_product_17(322) <= temp_mult_103(322);
partial_product_17(323) <= temp_mult_103(323);
partial_product_17(324) <= temp_mult_103(324);
partial_product_17(325) <= temp_mult_103(325);
partial_product_17(326) <= temp_mult_103(326);
partial_product_17(327) <= temp_mult_103(327);
partial_product_17(328) <= temp_mult_103(328);
partial_product_17(329) <= temp_mult_103(329);
partial_product_17(330) <= temp_mult_103(330);
partial_product_17(331) <= temp_mult_103(331);
partial_product_17(332) <= temp_mult_103(332);
partial_product_17(333) <= temp_mult_103(333);
partial_product_17(334) <= temp_mult_103(334);
partial_product_17(335) <= temp_mult_103(335);
partial_product_17(336) <= temp_mult_103(336);
partial_product_17(337) <= temp_mult_103(337);
partial_product_17(338) <= temp_mult_103(338);
partial_product_17(339) <= temp_mult_103(339);
partial_product_17(340) <= temp_mult_103(340);
partial_product_17(341) <= temp_mult_103(341);
partial_product_17(342) <= temp_mult_103(342);
partial_product_17(343) <= temp_mult_103(343);
partial_product_17(344) <= '0';
partial_product_17(345) <= '0';
partial_product_17(346) <= '0';
partial_product_17(347) <= '0';
partial_product_17(348) <= '0';
partial_product_17(349) <= '0';
partial_product_17(350) <= '0';
partial_product_17(351) <= '0';
partial_product_17(352) <= '0';
partial_product_17(353) <= '0';
partial_product_17(354) <= '0';
partial_product_17(355) <= '0';
partial_product_17(356) <= '0';
partial_product_17(357) <= '0';
partial_product_17(358) <= '0';
partial_product_17(359) <= '0';
partial_product_17(360) <= '0';
partial_product_17(361) <= '0';
partial_product_17(362) <= '0';
partial_product_17(363) <= '0';
partial_product_17(364) <= '0';
partial_product_17(365) <= '0';
partial_product_17(366) <= '0';
partial_product_17(367) <= '0';
partial_product_17(368) <= '0';
partial_product_17(369) <= '0';
partial_product_17(370) <= '0';
partial_product_17(371) <= '0';
partial_product_17(372) <= '0';
partial_product_17(373) <= '0';
partial_product_17(374) <= '0';
partial_product_17(375) <= '0';
partial_product_17(376) <= '0';
partial_product_17(377) <= '0';
partial_product_17(378) <= '0';
partial_product_17(379) <= '0';
partial_product_17(380) <= '0';
partial_product_17(381) <= '0';
partial_product_17(382) <= '0';
partial_product_17(383) <= '0';
partial_product_17(384) <= '0';
partial_product_17(385) <= '0';
partial_product_17(386) <= '0';
partial_product_17(387) <= '0';
partial_product_17(388) <= '0';
partial_product_17(389) <= '0';
partial_product_17(390) <= '0';
partial_product_17(391) <= '0';
partial_product_17(392) <= '0';
partial_product_17(393) <= '0';
partial_product_17(394) <= '0';
partial_product_17(395) <= '0';
partial_product_17(396) <= '0';
partial_product_17(397) <= '0';
partial_product_17(398) <= '0';
partial_product_17(399) <= '0';
partial_product_17(400) <= '0';
partial_product_17(401) <= '0';
partial_product_17(402) <= '0';
partial_product_17(403) <= '0';
partial_product_17(404) <= '0';
partial_product_17(405) <= '0';
partial_product_17(406) <= '0';
partial_product_17(407) <= '0';
partial_product_17(408) <= '0';
partial_product_17(409) <= '0';
partial_product_17(410) <= '0';
partial_product_17(411) <= '0';
partial_product_17(412) <= '0';
partial_product_17(413) <= '0';
partial_product_17(414) <= '0';
partial_product_17(415) <= '0';
partial_product_17(416) <= '0';
partial_product_17(417) <= '0';
partial_product_17(418) <= '0';
partial_product_17(419) <= '0';
partial_product_17(420) <= '0';
partial_product_17(421) <= '0';
partial_product_17(422) <= '0';
partial_product_17(423) <= '0';
partial_product_17(424) <= '0';
partial_product_17(425) <= '0';
partial_product_17(426) <= '0';
partial_product_17(427) <= '0';
partial_product_17(428) <= '0';
partial_product_17(429) <= '0';
partial_product_17(430) <= '0';
partial_product_17(431) <= '0';
partial_product_17(432) <= '0';
partial_product_17(433) <= '0';
partial_product_17(434) <= '0';
partial_product_17(435) <= '0';
partial_product_17(436) <= '0';
partial_product_17(437) <= '0';
partial_product_17(438) <= '0';
partial_product_17(439) <= '0';
partial_product_17(440) <= '0';
partial_product_17(441) <= '0';
partial_product_17(442) <= '0';
partial_product_17(443) <= '0';
partial_product_17(444) <= '0';
partial_product_17(445) <= '0';
partial_product_17(446) <= '0';
partial_product_17(447) <= '0';
partial_product_17(448) <= '0';
partial_product_17(449) <= '0';
partial_product_17(450) <= '0';
partial_product_17(451) <= '0';
partial_product_17(452) <= '0';
partial_product_17(453) <= '0';
partial_product_17(454) <= '0';
partial_product_17(455) <= '0';
partial_product_17(456) <= '0';
partial_product_17(457) <= '0';
partial_product_17(458) <= '0';
partial_product_17(459) <= '0';
partial_product_17(460) <= '0';
partial_product_17(461) <= '0';
partial_product_17(462) <= '0';
partial_product_17(463) <= '0';
partial_product_17(464) <= '0';
partial_product_17(465) <= '0';
partial_product_17(466) <= '0';
partial_product_17(467) <= '0';
partial_product_17(468) <= '0';
partial_product_17(469) <= '0';
partial_product_17(470) <= '0';
partial_product_17(471) <= '0';
partial_product_17(472) <= '0';
partial_product_17(473) <= '0';
partial_product_17(474) <= '0';
partial_product_17(475) <= '0';
partial_product_17(476) <= '0';
partial_product_17(477) <= '0';
partial_product_17(478) <= '0';
partial_product_17(479) <= '0';
partial_product_17(480) <= '0';
partial_product_17(481) <= '0';
partial_product_17(482) <= '0';
partial_product_17(483) <= '0';
partial_product_17(484) <= '0';
partial_product_17(485) <= '0';
partial_product_17(486) <= '0';
partial_product_17(487) <= '0';
partial_product_17(488) <= '0';
partial_product_17(489) <= '0';
partial_product_17(490) <= '0';
partial_product_17(491) <= '0';
partial_product_17(492) <= '0';
partial_product_17(493) <= '0';
partial_product_17(494) <= '0';
partial_product_17(495) <= '0';
partial_product_17(496) <= '0';
partial_product_17(497) <= '0';
partial_product_17(498) <= '0';
partial_product_17(499) <= '0';
partial_product_17(500) <= '0';
partial_product_17(501) <= '0';
partial_product_17(502) <= '0';
partial_product_17(503) <= '0';
partial_product_17(504) <= '0';
partial_product_17(505) <= '0';
partial_product_17(506) <= '0';
partial_product_17(507) <= '0';
partial_product_17(508) <= '0';
partial_product_17(509) <= '0';
partial_product_17(510) <= '0';
partial_product_17(511) <= '0';
partial_product_17(512) <= '0';
partial_product_18(0) <= '0';
partial_product_18(1) <= '0';
partial_product_18(2) <= '0';
partial_product_18(3) <= '0';
partial_product_18(4) <= '0';
partial_product_18(5) <= '0';
partial_product_18(6) <= '0';
partial_product_18(7) <= '0';
partial_product_18(8) <= '0';
partial_product_18(9) <= '0';
partial_product_18(10) <= '0';
partial_product_18(11) <= '0';
partial_product_18(12) <= '0';
partial_product_18(13) <= '0';
partial_product_18(14) <= '0';
partial_product_18(15) <= '0';
partial_product_18(16) <= '0';
partial_product_18(17) <= '0';
partial_product_18(18) <= '0';
partial_product_18(19) <= '0';
partial_product_18(20) <= '0';
partial_product_18(21) <= '0';
partial_product_18(22) <= '0';
partial_product_18(23) <= '0';
partial_product_18(24) <= '0';
partial_product_18(25) <= '0';
partial_product_18(26) <= '0';
partial_product_18(27) <= '0';
partial_product_18(28) <= '0';
partial_product_18(29) <= '0';
partial_product_18(30) <= '0';
partial_product_18(31) <= '0';
partial_product_18(32) <= '0';
partial_product_18(33) <= '0';
partial_product_18(34) <= '0';
partial_product_18(35) <= '0';
partial_product_18(36) <= '0';
partial_product_18(37) <= '0';
partial_product_18(38) <= '0';
partial_product_18(39) <= '0';
partial_product_18(40) <= '0';
partial_product_18(41) <= '0';
partial_product_18(42) <= '0';
partial_product_18(43) <= '0';
partial_product_18(44) <= '0';
partial_product_18(45) <= '0';
partial_product_18(46) <= '0';
partial_product_18(47) <= '0';
partial_product_18(48) <= '0';
partial_product_18(49) <= '0';
partial_product_18(50) <= '0';
partial_product_18(51) <= '0';
partial_product_18(52) <= '0';
partial_product_18(53) <= '0';
partial_product_18(54) <= '0';
partial_product_18(55) <= '0';
partial_product_18(56) <= '0';
partial_product_18(57) <= '0';
partial_product_18(58) <= '0';
partial_product_18(59) <= '0';
partial_product_18(60) <= '0';
partial_product_18(61) <= '0';
partial_product_18(62) <= '0';
partial_product_18(63) <= '0';
partial_product_18(64) <= '0';
partial_product_18(65) <= '0';
partial_product_18(66) <= '0';
partial_product_18(67) <= '0';
partial_product_18(68) <= '0';
partial_product_18(69) <= '0';
partial_product_18(70) <= '0';
partial_product_18(71) <= '0';
partial_product_18(72) <= '0';
partial_product_18(73) <= '0';
partial_product_18(74) <= '0';
partial_product_18(75) <= '0';
partial_product_18(76) <= '0';
partial_product_18(77) <= '0';
partial_product_18(78) <= '0';
partial_product_18(79) <= '0';
partial_product_18(80) <= '0';
partial_product_18(81) <= '0';
partial_product_18(82) <= '0';
partial_product_18(83) <= '0';
partial_product_18(84) <= '0';
partial_product_18(85) <= '0';
partial_product_18(86) <= '0';
partial_product_18(87) <= '0';
partial_product_18(88) <= '0';
partial_product_18(89) <= '0';
partial_product_18(90) <= '0';
partial_product_18(91) <= '0';
partial_product_18(92) <= '0';
partial_product_18(93) <= '0';
partial_product_18(94) <= '0';
partial_product_18(95) <= '0';
partial_product_18(96) <= '0';
partial_product_18(97) <= '0';
partial_product_18(98) <= '0';
partial_product_18(99) <= '0';
partial_product_18(100) <= '0';
partial_product_18(101) <= '0';
partial_product_18(102) <= '0';
partial_product_18(103) <= '0';
partial_product_18(104) <= '0';
partial_product_18(105) <= '0';
partial_product_18(106) <= '0';
partial_product_18(107) <= '0';
partial_product_18(108) <= '0';
partial_product_18(109) <= '0';
partial_product_18(110) <= '0';
partial_product_18(111) <= '0';
partial_product_18(112) <= '0';
partial_product_18(113) <= '0';
partial_product_18(114) <= '0';
partial_product_18(115) <= '0';
partial_product_18(116) <= '0';
partial_product_18(117) <= '0';
partial_product_18(118) <= '0';
partial_product_18(119) <= '0';
partial_product_18(120) <= '0';
partial_product_18(121) <= '0';
partial_product_18(122) <= '0';
partial_product_18(123) <= '0';
partial_product_18(124) <= '0';
partial_product_18(125) <= '0';
partial_product_18(126) <= '0';
partial_product_18(127) <= '0';
partial_product_18(128) <= '0';
partial_product_18(129) <= '0';
partial_product_18(130) <= '0';
partial_product_18(131) <= '0';
partial_product_18(132) <= '0';
partial_product_18(133) <= '0';
partial_product_18(134) <= '0';
partial_product_18(135) <= '0';
partial_product_18(136) <= '0';
partial_product_18(137) <= '0';
partial_product_18(138) <= '0';
partial_product_18(139) <= '0';
partial_product_18(140) <= '0';
partial_product_18(141) <= '0';
partial_product_18(142) <= '0';
partial_product_18(143) <= '0';
partial_product_18(144) <= '0';
partial_product_18(145) <= '0';
partial_product_18(146) <= '0';
partial_product_18(147) <= '0';
partial_product_18(148) <= '0';
partial_product_18(149) <= '0';
partial_product_18(150) <= '0';
partial_product_18(151) <= '0';
partial_product_18(152) <= '0';
partial_product_18(153) <= '0';
partial_product_18(154) <= '0';
partial_product_18(155) <= '0';
partial_product_18(156) <= '0';
partial_product_18(157) <= '0';
partial_product_18(158) <= '0';
partial_product_18(159) <= '0';
partial_product_18(160) <= '0';
partial_product_18(161) <= '0';
partial_product_18(162) <= '0';
partial_product_18(163) <= '0';
partial_product_18(164) <= '0';
partial_product_18(165) <= '0';
partial_product_18(166) <= '0';
partial_product_18(167) <= '0';
partial_product_18(168) <= '0';
partial_product_18(169) <= '0';
partial_product_18(170) <= '0';
partial_product_18(171) <= '0';
partial_product_18(172) <= '0';
partial_product_18(173) <= '0';
partial_product_18(174) <= '0';
partial_product_18(175) <= '0';
partial_product_18(176) <= '0';
partial_product_18(177) <= '0';
partial_product_18(178) <= '0';
partial_product_18(179) <= '0';
partial_product_18(180) <= '0';
partial_product_18(181) <= '0';
partial_product_18(182) <= '0';
partial_product_18(183) <= '0';
partial_product_18(184) <= '0';
partial_product_18(185) <= '0';
partial_product_18(186) <= '0';
partial_product_18(187) <= temp_mult_83(187);
partial_product_18(188) <= temp_mult_83(188);
partial_product_18(189) <= temp_mult_83(189);
partial_product_18(190) <= temp_mult_83(190);
partial_product_18(191) <= temp_mult_83(191);
partial_product_18(192) <= temp_mult_83(192);
partial_product_18(193) <= temp_mult_83(193);
partial_product_18(194) <= temp_mult_83(194);
partial_product_18(195) <= temp_mult_83(195);
partial_product_18(196) <= temp_mult_83(196);
partial_product_18(197) <= temp_mult_83(197);
partial_product_18(198) <= temp_mult_83(198);
partial_product_18(199) <= temp_mult_83(199);
partial_product_18(200) <= temp_mult_83(200);
partial_product_18(201) <= temp_mult_83(201);
partial_product_18(202) <= temp_mult_83(202);
partial_product_18(203) <= temp_mult_83(203);
partial_product_18(204) <= temp_mult_83(204);
partial_product_18(205) <= temp_mult_83(205);
partial_product_18(206) <= temp_mult_83(206);
partial_product_18(207) <= temp_mult_83(207);
partial_product_18(208) <= temp_mult_83(208);
partial_product_18(209) <= temp_mult_83(209);
partial_product_18(210) <= temp_mult_83(210);
partial_product_18(211) <= temp_mult_83(211);
partial_product_18(212) <= temp_mult_83(212);
partial_product_18(213) <= temp_mult_83(213);
partial_product_18(214) <= temp_mult_83(214);
partial_product_18(215) <= temp_mult_83(215);
partial_product_18(216) <= temp_mult_83(216);
partial_product_18(217) <= temp_mult_83(217);
partial_product_18(218) <= temp_mult_83(218);
partial_product_18(219) <= temp_mult_83(219);
partial_product_18(220) <= temp_mult_83(220);
partial_product_18(221) <= temp_mult_83(221);
partial_product_18(222) <= temp_mult_83(222);
partial_product_18(223) <= temp_mult_83(223);
partial_product_18(224) <= temp_mult_83(224);
partial_product_18(225) <= temp_mult_83(225);
partial_product_18(226) <= temp_mult_83(226);
partial_product_18(227) <= temp_mult_83(227);
partial_product_18(228) <= temp_mult_92(228);
partial_product_18(229) <= temp_mult_92(229);
partial_product_18(230) <= temp_mult_92(230);
partial_product_18(231) <= temp_mult_92(231);
partial_product_18(232) <= temp_mult_92(232);
partial_product_18(233) <= temp_mult_92(233);
partial_product_18(234) <= temp_mult_92(234);
partial_product_18(235) <= temp_mult_92(235);
partial_product_18(236) <= temp_mult_92(236);
partial_product_18(237) <= temp_mult_92(237);
partial_product_18(238) <= temp_mult_92(238);
partial_product_18(239) <= temp_mult_92(239);
partial_product_18(240) <= temp_mult_92(240);
partial_product_18(241) <= temp_mult_92(241);
partial_product_18(242) <= temp_mult_92(242);
partial_product_18(243) <= temp_mult_92(243);
partial_product_18(244) <= temp_mult_92(244);
partial_product_18(245) <= temp_mult_92(245);
partial_product_18(246) <= temp_mult_92(246);
partial_product_18(247) <= temp_mult_92(247);
partial_product_18(248) <= temp_mult_92(248);
partial_product_18(249) <= temp_mult_92(249);
partial_product_18(250) <= temp_mult_92(250);
partial_product_18(251) <= temp_mult_92(251);
partial_product_18(252) <= temp_mult_92(252);
partial_product_18(253) <= temp_mult_92(253);
partial_product_18(254) <= temp_mult_92(254);
partial_product_18(255) <= temp_mult_92(255);
partial_product_18(256) <= temp_mult_92(256);
partial_product_18(257) <= temp_mult_92(257);
partial_product_18(258) <= temp_mult_92(258);
partial_product_18(259) <= temp_mult_92(259);
partial_product_18(260) <= temp_mult_92(260);
partial_product_18(261) <= temp_mult_92(261);
partial_product_18(262) <= temp_mult_92(262);
partial_product_18(263) <= temp_mult_92(263);
partial_product_18(264) <= temp_mult_92(264);
partial_product_18(265) <= temp_mult_92(265);
partial_product_18(266) <= temp_mult_92(266);
partial_product_18(267) <= temp_mult_92(267);
partial_product_18(268) <= temp_mult_92(268);
partial_product_18(269) <= temp_mult_101(269);
partial_product_18(270) <= temp_mult_101(270);
partial_product_18(271) <= temp_mult_101(271);
partial_product_18(272) <= temp_mult_101(272);
partial_product_18(273) <= temp_mult_101(273);
partial_product_18(274) <= temp_mult_101(274);
partial_product_18(275) <= temp_mult_101(275);
partial_product_18(276) <= temp_mult_101(276);
partial_product_18(277) <= temp_mult_101(277);
partial_product_18(278) <= temp_mult_101(278);
partial_product_18(279) <= temp_mult_101(279);
partial_product_18(280) <= temp_mult_101(280);
partial_product_18(281) <= temp_mult_101(281);
partial_product_18(282) <= temp_mult_101(282);
partial_product_18(283) <= temp_mult_101(283);
partial_product_18(284) <= temp_mult_101(284);
partial_product_18(285) <= temp_mult_101(285);
partial_product_18(286) <= temp_mult_101(286);
partial_product_18(287) <= temp_mult_101(287);
partial_product_18(288) <= temp_mult_101(288);
partial_product_18(289) <= temp_mult_101(289);
partial_product_18(290) <= temp_mult_101(290);
partial_product_18(291) <= temp_mult_101(291);
partial_product_18(292) <= temp_mult_101(292);
partial_product_18(293) <= temp_mult_101(293);
partial_product_18(294) <= temp_mult_101(294);
partial_product_18(295) <= temp_mult_101(295);
partial_product_18(296) <= temp_mult_101(296);
partial_product_18(297) <= temp_mult_101(297);
partial_product_18(298) <= temp_mult_101(298);
partial_product_18(299) <= temp_mult_101(299);
partial_product_18(300) <= temp_mult_101(300);
partial_product_18(301) <= temp_mult_101(301);
partial_product_18(302) <= temp_mult_101(302);
partial_product_18(303) <= temp_mult_101(303);
partial_product_18(304) <= temp_mult_101(304);
partial_product_18(305) <= temp_mult_101(305);
partial_product_18(306) <= temp_mult_101(306);
partial_product_18(307) <= temp_mult_101(307);
partial_product_18(308) <= temp_mult_101(308);
partial_product_18(309) <= temp_mult_101(309);
partial_product_18(310) <= '0';
partial_product_18(311) <= '0';
partial_product_18(312) <= '0';
partial_product_18(313) <= '0';
partial_product_18(314) <= '0';
partial_product_18(315) <= '0';
partial_product_18(316) <= '0';
partial_product_18(317) <= '0';
partial_product_18(318) <= '0';
partial_product_18(319) <= '0';
partial_product_18(320) <= '0';
partial_product_18(321) <= '0';
partial_product_18(322) <= '0';
partial_product_18(323) <= '0';
partial_product_18(324) <= '0';
partial_product_18(325) <= '0';
partial_product_18(326) <= '0';
partial_product_18(327) <= '0';
partial_product_18(328) <= '0';
partial_product_18(329) <= '0';
partial_product_18(330) <= '0';
partial_product_18(331) <= '0';
partial_product_18(332) <= '0';
partial_product_18(333) <= '0';
partial_product_18(334) <= '0';
partial_product_18(335) <= '0';
partial_product_18(336) <= '0';
partial_product_18(337) <= '0';
partial_product_18(338) <= '0';
partial_product_18(339) <= '0';
partial_product_18(340) <= '0';
partial_product_18(341) <= '0';
partial_product_18(342) <= '0';
partial_product_18(343) <= '0';
partial_product_18(344) <= '0';
partial_product_18(345) <= '0';
partial_product_18(346) <= '0';
partial_product_18(347) <= '0';
partial_product_18(348) <= '0';
partial_product_18(349) <= '0';
partial_product_18(350) <= '0';
partial_product_18(351) <= '0';
partial_product_18(352) <= '0';
partial_product_18(353) <= '0';
partial_product_18(354) <= '0';
partial_product_18(355) <= '0';
partial_product_18(356) <= '0';
partial_product_18(357) <= '0';
partial_product_18(358) <= '0';
partial_product_18(359) <= '0';
partial_product_18(360) <= '0';
partial_product_18(361) <= '0';
partial_product_18(362) <= '0';
partial_product_18(363) <= '0';
partial_product_18(364) <= '0';
partial_product_18(365) <= '0';
partial_product_18(366) <= '0';
partial_product_18(367) <= '0';
partial_product_18(368) <= '0';
partial_product_18(369) <= '0';
partial_product_18(370) <= '0';
partial_product_18(371) <= '0';
partial_product_18(372) <= '0';
partial_product_18(373) <= '0';
partial_product_18(374) <= '0';
partial_product_18(375) <= '0';
partial_product_18(376) <= '0';
partial_product_18(377) <= '0';
partial_product_18(378) <= '0';
partial_product_18(379) <= '0';
partial_product_18(380) <= '0';
partial_product_18(381) <= '0';
partial_product_18(382) <= '0';
partial_product_18(383) <= '0';
partial_product_18(384) <= '0';
partial_product_18(385) <= '0';
partial_product_18(386) <= '0';
partial_product_18(387) <= '0';
partial_product_18(388) <= '0';
partial_product_18(389) <= '0';
partial_product_18(390) <= '0';
partial_product_18(391) <= '0';
partial_product_18(392) <= '0';
partial_product_18(393) <= '0';
partial_product_18(394) <= '0';
partial_product_18(395) <= '0';
partial_product_18(396) <= '0';
partial_product_18(397) <= '0';
partial_product_18(398) <= '0';
partial_product_18(399) <= '0';
partial_product_18(400) <= '0';
partial_product_18(401) <= '0';
partial_product_18(402) <= '0';
partial_product_18(403) <= '0';
partial_product_18(404) <= '0';
partial_product_18(405) <= '0';
partial_product_18(406) <= '0';
partial_product_18(407) <= '0';
partial_product_18(408) <= '0';
partial_product_18(409) <= '0';
partial_product_18(410) <= '0';
partial_product_18(411) <= '0';
partial_product_18(412) <= '0';
partial_product_18(413) <= '0';
partial_product_18(414) <= '0';
partial_product_18(415) <= '0';
partial_product_18(416) <= '0';
partial_product_18(417) <= '0';
partial_product_18(418) <= '0';
partial_product_18(419) <= '0';
partial_product_18(420) <= '0';
partial_product_18(421) <= '0';
partial_product_18(422) <= '0';
partial_product_18(423) <= '0';
partial_product_18(424) <= '0';
partial_product_18(425) <= '0';
partial_product_18(426) <= '0';
partial_product_18(427) <= '0';
partial_product_18(428) <= '0';
partial_product_18(429) <= '0';
partial_product_18(430) <= '0';
partial_product_18(431) <= '0';
partial_product_18(432) <= '0';
partial_product_18(433) <= '0';
partial_product_18(434) <= '0';
partial_product_18(435) <= '0';
partial_product_18(436) <= '0';
partial_product_18(437) <= '0';
partial_product_18(438) <= '0';
partial_product_18(439) <= '0';
partial_product_18(440) <= '0';
partial_product_18(441) <= '0';
partial_product_18(442) <= '0';
partial_product_18(443) <= '0';
partial_product_18(444) <= '0';
partial_product_18(445) <= '0';
partial_product_18(446) <= '0';
partial_product_18(447) <= '0';
partial_product_18(448) <= '0';
partial_product_18(449) <= '0';
partial_product_18(450) <= '0';
partial_product_18(451) <= '0';
partial_product_18(452) <= '0';
partial_product_18(453) <= '0';
partial_product_18(454) <= '0';
partial_product_18(455) <= '0';
partial_product_18(456) <= '0';
partial_product_18(457) <= '0';
partial_product_18(458) <= '0';
partial_product_18(459) <= '0';
partial_product_18(460) <= '0';
partial_product_18(461) <= '0';
partial_product_18(462) <= '0';
partial_product_18(463) <= '0';
partial_product_18(464) <= '0';
partial_product_18(465) <= '0';
partial_product_18(466) <= '0';
partial_product_18(467) <= '0';
partial_product_18(468) <= '0';
partial_product_18(469) <= '0';
partial_product_18(470) <= '0';
partial_product_18(471) <= '0';
partial_product_18(472) <= '0';
partial_product_18(473) <= '0';
partial_product_18(474) <= '0';
partial_product_18(475) <= '0';
partial_product_18(476) <= '0';
partial_product_18(477) <= '0';
partial_product_18(478) <= '0';
partial_product_18(479) <= '0';
partial_product_18(480) <= '0';
partial_product_18(481) <= '0';
partial_product_18(482) <= '0';
partial_product_18(483) <= '0';
partial_product_18(484) <= '0';
partial_product_18(485) <= '0';
partial_product_18(486) <= '0';
partial_product_18(487) <= '0';
partial_product_18(488) <= '0';
partial_product_18(489) <= '0';
partial_product_18(490) <= '0';
partial_product_18(491) <= '0';
partial_product_18(492) <= '0';
partial_product_18(493) <= '0';
partial_product_18(494) <= '0';
partial_product_18(495) <= '0';
partial_product_18(496) <= '0';
partial_product_18(497) <= '0';
partial_product_18(498) <= '0';
partial_product_18(499) <= '0';
partial_product_18(500) <= '0';
partial_product_18(501) <= '0';
partial_product_18(502) <= '0';
partial_product_18(503) <= '0';
partial_product_18(504) <= '0';
partial_product_18(505) <= '0';
partial_product_18(506) <= '0';
partial_product_18(507) <= '0';
partial_product_18(508) <= '0';
partial_product_18(509) <= '0';
partial_product_18(510) <= '0';
partial_product_18(511) <= '0';
partial_product_18(512) <= '0';
partial_product_19(0) <= '0';
partial_product_19(1) <= '0';
partial_product_19(2) <= '0';
partial_product_19(3) <= '0';
partial_product_19(4) <= '0';
partial_product_19(5) <= '0';
partial_product_19(6) <= '0';
partial_product_19(7) <= '0';
partial_product_19(8) <= '0';
partial_product_19(9) <= '0';
partial_product_19(10) <= '0';
partial_product_19(11) <= '0';
partial_product_19(12) <= '0';
partial_product_19(13) <= '0';
partial_product_19(14) <= '0';
partial_product_19(15) <= '0';
partial_product_19(16) <= '0';
partial_product_19(17) <= '0';
partial_product_19(18) <= '0';
partial_product_19(19) <= '0';
partial_product_19(20) <= '0';
partial_product_19(21) <= '0';
partial_product_19(22) <= '0';
partial_product_19(23) <= '0';
partial_product_19(24) <= '0';
partial_product_19(25) <= '0';
partial_product_19(26) <= '0';
partial_product_19(27) <= '0';
partial_product_19(28) <= '0';
partial_product_19(29) <= '0';
partial_product_19(30) <= '0';
partial_product_19(31) <= '0';
partial_product_19(32) <= '0';
partial_product_19(33) <= '0';
partial_product_19(34) <= '0';
partial_product_19(35) <= '0';
partial_product_19(36) <= '0';
partial_product_19(37) <= '0';
partial_product_19(38) <= '0';
partial_product_19(39) <= '0';
partial_product_19(40) <= '0';
partial_product_19(41) <= '0';
partial_product_19(42) <= '0';
partial_product_19(43) <= '0';
partial_product_19(44) <= '0';
partial_product_19(45) <= '0';
partial_product_19(46) <= '0';
partial_product_19(47) <= '0';
partial_product_19(48) <= '0';
partial_product_19(49) <= '0';
partial_product_19(50) <= '0';
partial_product_19(51) <= '0';
partial_product_19(52) <= '0';
partial_product_19(53) <= '0';
partial_product_19(54) <= '0';
partial_product_19(55) <= '0';
partial_product_19(56) <= '0';
partial_product_19(57) <= '0';
partial_product_19(58) <= '0';
partial_product_19(59) <= '0';
partial_product_19(60) <= '0';
partial_product_19(61) <= '0';
partial_product_19(62) <= '0';
partial_product_19(63) <= '0';
partial_product_19(64) <= '0';
partial_product_19(65) <= '0';
partial_product_19(66) <= '0';
partial_product_19(67) <= '0';
partial_product_19(68) <= '0';
partial_product_19(69) <= '0';
partial_product_19(70) <= '0';
partial_product_19(71) <= '0';
partial_product_19(72) <= '0';
partial_product_19(73) <= '0';
partial_product_19(74) <= '0';
partial_product_19(75) <= '0';
partial_product_19(76) <= '0';
partial_product_19(77) <= '0';
partial_product_19(78) <= '0';
partial_product_19(79) <= '0';
partial_product_19(80) <= '0';
partial_product_19(81) <= '0';
partial_product_19(82) <= '0';
partial_product_19(83) <= '0';
partial_product_19(84) <= '0';
partial_product_19(85) <= '0';
partial_product_19(86) <= '0';
partial_product_19(87) <= '0';
partial_product_19(88) <= '0';
partial_product_19(89) <= '0';
partial_product_19(90) <= '0';
partial_product_19(91) <= '0';
partial_product_19(92) <= '0';
partial_product_19(93) <= '0';
partial_product_19(94) <= '0';
partial_product_19(95) <= '0';
partial_product_19(96) <= '0';
partial_product_19(97) <= '0';
partial_product_19(98) <= '0';
partial_product_19(99) <= '0';
partial_product_19(100) <= '0';
partial_product_19(101) <= '0';
partial_product_19(102) <= '0';
partial_product_19(103) <= '0';
partial_product_19(104) <= '0';
partial_product_19(105) <= '0';
partial_product_19(106) <= '0';
partial_product_19(107) <= '0';
partial_product_19(108) <= '0';
partial_product_19(109) <= '0';
partial_product_19(110) <= '0';
partial_product_19(111) <= '0';
partial_product_19(112) <= '0';
partial_product_19(113) <= '0';
partial_product_19(114) <= '0';
partial_product_19(115) <= '0';
partial_product_19(116) <= '0';
partial_product_19(117) <= '0';
partial_product_19(118) <= '0';
partial_product_19(119) <= '0';
partial_product_19(120) <= '0';
partial_product_19(121) <= '0';
partial_product_19(122) <= '0';
partial_product_19(123) <= '0';
partial_product_19(124) <= '0';
partial_product_19(125) <= '0';
partial_product_19(126) <= '0';
partial_product_19(127) <= '0';
partial_product_19(128) <= '0';
partial_product_19(129) <= '0';
partial_product_19(130) <= '0';
partial_product_19(131) <= '0';
partial_product_19(132) <= '0';
partial_product_19(133) <= '0';
partial_product_19(134) <= '0';
partial_product_19(135) <= '0';
partial_product_19(136) <= '0';
partial_product_19(137) <= '0';
partial_product_19(138) <= '0';
partial_product_19(139) <= '0';
partial_product_19(140) <= '0';
partial_product_19(141) <= '0';
partial_product_19(142) <= '0';
partial_product_19(143) <= '0';
partial_product_19(144) <= '0';
partial_product_19(145) <= '0';
partial_product_19(146) <= '0';
partial_product_19(147) <= '0';
partial_product_19(148) <= '0';
partial_product_19(149) <= '0';
partial_product_19(150) <= '0';
partial_product_19(151) <= '0';
partial_product_19(152) <= '0';
partial_product_19(153) <= '0';
partial_product_19(154) <= '0';
partial_product_19(155) <= '0';
partial_product_19(156) <= '0';
partial_product_19(157) <= '0';
partial_product_19(158) <= '0';
partial_product_19(159) <= '0';
partial_product_19(160) <= '0';
partial_product_19(161) <= '0';
partial_product_19(162) <= '0';
partial_product_19(163) <= '0';
partial_product_19(164) <= '0';
partial_product_19(165) <= '0';
partial_product_19(166) <= '0';
partial_product_19(167) <= '0';
partial_product_19(168) <= '0';
partial_product_19(169) <= '0';
partial_product_19(170) <= '0';
partial_product_19(171) <= '0';
partial_product_19(172) <= '0';
partial_product_19(173) <= '0';
partial_product_19(174) <= '0';
partial_product_19(175) <= '0';
partial_product_19(176) <= '0';
partial_product_19(177) <= '0';
partial_product_19(178) <= '0';
partial_product_19(179) <= '0';
partial_product_19(180) <= '0';
partial_product_19(181) <= '0';
partial_product_19(182) <= '0';
partial_product_19(183) <= '0';
partial_product_19(184) <= '0';
partial_product_19(185) <= '0';
partial_product_19(186) <= '0';
partial_product_19(187) <= '0';
partial_product_19(188) <= '0';
partial_product_19(189) <= '0';
partial_product_19(190) <= '0';
partial_product_19(191) <= '0';
partial_product_19(192) <= temp_mult_64(192);
partial_product_19(193) <= temp_mult_64(193);
partial_product_19(194) <= temp_mult_64(194);
partial_product_19(195) <= temp_mult_64(195);
partial_product_19(196) <= temp_mult_64(196);
partial_product_19(197) <= temp_mult_64(197);
partial_product_19(198) <= temp_mult_64(198);
partial_product_19(199) <= temp_mult_64(199);
partial_product_19(200) <= temp_mult_64(200);
partial_product_19(201) <= temp_mult_64(201);
partial_product_19(202) <= temp_mult_64(202);
partial_product_19(203) <= temp_mult_64(203);
partial_product_19(204) <= temp_mult_64(204);
partial_product_19(205) <= temp_mult_64(205);
partial_product_19(206) <= temp_mult_64(206);
partial_product_19(207) <= temp_mult_64(207);
partial_product_19(208) <= temp_mult_64(208);
partial_product_19(209) <= temp_mult_64(209);
partial_product_19(210) <= temp_mult_64(210);
partial_product_19(211) <= temp_mult_64(211);
partial_product_19(212) <= temp_mult_64(212);
partial_product_19(213) <= temp_mult_64(213);
partial_product_19(214) <= temp_mult_64(214);
partial_product_19(215) <= temp_mult_64(215);
partial_product_19(216) <= temp_mult_64(216);
partial_product_19(217) <= temp_mult_64(217);
partial_product_19(218) <= temp_mult_64(218);
partial_product_19(219) <= temp_mult_64(219);
partial_product_19(220) <= temp_mult_64(220);
partial_product_19(221) <= temp_mult_64(221);
partial_product_19(222) <= temp_mult_64(222);
partial_product_19(223) <= temp_mult_64(223);
partial_product_19(224) <= temp_mult_64(224);
partial_product_19(225) <= temp_mult_64(225);
partial_product_19(226) <= temp_mult_64(226);
partial_product_19(227) <= temp_mult_64(227);
partial_product_19(228) <= temp_mult_64(228);
partial_product_19(229) <= temp_mult_64(229);
partial_product_19(230) <= temp_mult_64(230);
partial_product_19(231) <= temp_mult_64(231);
partial_product_19(232) <= temp_mult_64(232);
partial_product_19(233) <= temp_mult_73(233);
partial_product_19(234) <= temp_mult_73(234);
partial_product_19(235) <= temp_mult_73(235);
partial_product_19(236) <= temp_mult_73(236);
partial_product_19(237) <= temp_mult_73(237);
partial_product_19(238) <= temp_mult_73(238);
partial_product_19(239) <= temp_mult_73(239);
partial_product_19(240) <= temp_mult_73(240);
partial_product_19(241) <= temp_mult_73(241);
partial_product_19(242) <= temp_mult_73(242);
partial_product_19(243) <= temp_mult_73(243);
partial_product_19(244) <= temp_mult_73(244);
partial_product_19(245) <= temp_mult_73(245);
partial_product_19(246) <= temp_mult_73(246);
partial_product_19(247) <= temp_mult_73(247);
partial_product_19(248) <= temp_mult_73(248);
partial_product_19(249) <= temp_mult_73(249);
partial_product_19(250) <= temp_mult_73(250);
partial_product_19(251) <= temp_mult_73(251);
partial_product_19(252) <= temp_mult_73(252);
partial_product_19(253) <= temp_mult_73(253);
partial_product_19(254) <= temp_mult_73(254);
partial_product_19(255) <= temp_mult_73(255);
partial_product_19(256) <= temp_mult_73(256);
partial_product_19(257) <= temp_mult_73(257);
partial_product_19(258) <= temp_mult_73(258);
partial_product_19(259) <= temp_mult_73(259);
partial_product_19(260) <= temp_mult_73(260);
partial_product_19(261) <= temp_mult_73(261);
partial_product_19(262) <= temp_mult_73(262);
partial_product_19(263) <= temp_mult_73(263);
partial_product_19(264) <= temp_mult_73(264);
partial_product_19(265) <= temp_mult_73(265);
partial_product_19(266) <= temp_mult_73(266);
partial_product_19(267) <= temp_mult_73(267);
partial_product_19(268) <= temp_mult_73(268);
partial_product_19(269) <= temp_mult_73(269);
partial_product_19(270) <= temp_mult_73(270);
partial_product_19(271) <= temp_mult_73(271);
partial_product_19(272) <= temp_mult_73(272);
partial_product_19(273) <= temp_mult_73(273);
partial_product_19(274) <= '0';
partial_product_19(275) <= '0';
partial_product_19(276) <= '0';
partial_product_19(277) <= '0';
partial_product_19(278) <= '0';
partial_product_19(279) <= temp_mult_95(279);
partial_product_19(280) <= temp_mult_95(280);
partial_product_19(281) <= temp_mult_95(281);
partial_product_19(282) <= temp_mult_95(282);
partial_product_19(283) <= temp_mult_95(283);
partial_product_19(284) <= temp_mult_95(284);
partial_product_19(285) <= temp_mult_95(285);
partial_product_19(286) <= temp_mult_95(286);
partial_product_19(287) <= temp_mult_95(287);
partial_product_19(288) <= temp_mult_95(288);
partial_product_19(289) <= temp_mult_95(289);
partial_product_19(290) <= temp_mult_95(290);
partial_product_19(291) <= temp_mult_95(291);
partial_product_19(292) <= temp_mult_95(292);
partial_product_19(293) <= temp_mult_95(293);
partial_product_19(294) <= temp_mult_95(294);
partial_product_19(295) <= temp_mult_95(295);
partial_product_19(296) <= temp_mult_95(296);
partial_product_19(297) <= temp_mult_95(297);
partial_product_19(298) <= temp_mult_95(298);
partial_product_19(299) <= temp_mult_95(299);
partial_product_19(300) <= temp_mult_95(300);
partial_product_19(301) <= temp_mult_95(301);
partial_product_19(302) <= temp_mult_95(302);
partial_product_19(303) <= temp_mult_95(303);
partial_product_19(304) <= temp_mult_95(304);
partial_product_19(305) <= temp_mult_95(305);
partial_product_19(306) <= temp_mult_95(306);
partial_product_19(307) <= temp_mult_95(307);
partial_product_19(308) <= temp_mult_95(308);
partial_product_19(309) <= temp_mult_95(309);
partial_product_19(310) <= temp_mult_95(310);
partial_product_19(311) <= temp_mult_95(311);
partial_product_19(312) <= temp_mult_95(312);
partial_product_19(313) <= temp_mult_95(313);
partial_product_19(314) <= temp_mult_95(314);
partial_product_19(315) <= temp_mult_95(315);
partial_product_19(316) <= temp_mult_95(316);
partial_product_19(317) <= temp_mult_95(317);
partial_product_19(318) <= temp_mult_95(318);
partial_product_19(319) <= temp_mult_95(319);
partial_product_19(320) <= '0';
partial_product_19(321) <= '0';
partial_product_19(322) <= '0';
partial_product_19(323) <= '0';
partial_product_19(324) <= '0';
partial_product_19(325) <= '0';
partial_product_19(326) <= '0';
partial_product_19(327) <= '0';
partial_product_19(328) <= '0';
partial_product_19(329) <= '0';
partial_product_19(330) <= '0';
partial_product_19(331) <= '0';
partial_product_19(332) <= '0';
partial_product_19(333) <= '0';
partial_product_19(334) <= '0';
partial_product_19(335) <= '0';
partial_product_19(336) <= '0';
partial_product_19(337) <= '0';
partial_product_19(338) <= '0';
partial_product_19(339) <= '0';
partial_product_19(340) <= '0';
partial_product_19(341) <= '0';
partial_product_19(342) <= '0';
partial_product_19(343) <= '0';
partial_product_19(344) <= '0';
partial_product_19(345) <= '0';
partial_product_19(346) <= '0';
partial_product_19(347) <= '0';
partial_product_19(348) <= '0';
partial_product_19(349) <= '0';
partial_product_19(350) <= '0';
partial_product_19(351) <= '0';
partial_product_19(352) <= '0';
partial_product_19(353) <= '0';
partial_product_19(354) <= '0';
partial_product_19(355) <= '0';
partial_product_19(356) <= '0';
partial_product_19(357) <= '0';
partial_product_19(358) <= '0';
partial_product_19(359) <= '0';
partial_product_19(360) <= '0';
partial_product_19(361) <= '0';
partial_product_19(362) <= '0';
partial_product_19(363) <= '0';
partial_product_19(364) <= '0';
partial_product_19(365) <= '0';
partial_product_19(366) <= '0';
partial_product_19(367) <= '0';
partial_product_19(368) <= '0';
partial_product_19(369) <= '0';
partial_product_19(370) <= '0';
partial_product_19(371) <= '0';
partial_product_19(372) <= '0';
partial_product_19(373) <= '0';
partial_product_19(374) <= '0';
partial_product_19(375) <= '0';
partial_product_19(376) <= '0';
partial_product_19(377) <= '0';
partial_product_19(378) <= '0';
partial_product_19(379) <= '0';
partial_product_19(380) <= '0';
partial_product_19(381) <= '0';
partial_product_19(382) <= '0';
partial_product_19(383) <= '0';
partial_product_19(384) <= '0';
partial_product_19(385) <= '0';
partial_product_19(386) <= '0';
partial_product_19(387) <= '0';
partial_product_19(388) <= '0';
partial_product_19(389) <= '0';
partial_product_19(390) <= '0';
partial_product_19(391) <= '0';
partial_product_19(392) <= '0';
partial_product_19(393) <= '0';
partial_product_19(394) <= '0';
partial_product_19(395) <= '0';
partial_product_19(396) <= '0';
partial_product_19(397) <= '0';
partial_product_19(398) <= '0';
partial_product_19(399) <= '0';
partial_product_19(400) <= '0';
partial_product_19(401) <= '0';
partial_product_19(402) <= '0';
partial_product_19(403) <= '0';
partial_product_19(404) <= '0';
partial_product_19(405) <= '0';
partial_product_19(406) <= '0';
partial_product_19(407) <= '0';
partial_product_19(408) <= '0';
partial_product_19(409) <= '0';
partial_product_19(410) <= '0';
partial_product_19(411) <= '0';
partial_product_19(412) <= '0';
partial_product_19(413) <= '0';
partial_product_19(414) <= '0';
partial_product_19(415) <= '0';
partial_product_19(416) <= '0';
partial_product_19(417) <= '0';
partial_product_19(418) <= '0';
partial_product_19(419) <= '0';
partial_product_19(420) <= '0';
partial_product_19(421) <= '0';
partial_product_19(422) <= '0';
partial_product_19(423) <= '0';
partial_product_19(424) <= '0';
partial_product_19(425) <= '0';
partial_product_19(426) <= '0';
partial_product_19(427) <= '0';
partial_product_19(428) <= '0';
partial_product_19(429) <= '0';
partial_product_19(430) <= '0';
partial_product_19(431) <= '0';
partial_product_19(432) <= '0';
partial_product_19(433) <= '0';
partial_product_19(434) <= '0';
partial_product_19(435) <= '0';
partial_product_19(436) <= '0';
partial_product_19(437) <= '0';
partial_product_19(438) <= '0';
partial_product_19(439) <= '0';
partial_product_19(440) <= '0';
partial_product_19(441) <= '0';
partial_product_19(442) <= '0';
partial_product_19(443) <= '0';
partial_product_19(444) <= '0';
partial_product_19(445) <= '0';
partial_product_19(446) <= '0';
partial_product_19(447) <= '0';
partial_product_19(448) <= '0';
partial_product_19(449) <= '0';
partial_product_19(450) <= '0';
partial_product_19(451) <= '0';
partial_product_19(452) <= '0';
partial_product_19(453) <= '0';
partial_product_19(454) <= '0';
partial_product_19(455) <= '0';
partial_product_19(456) <= '0';
partial_product_19(457) <= '0';
partial_product_19(458) <= '0';
partial_product_19(459) <= '0';
partial_product_19(460) <= '0';
partial_product_19(461) <= '0';
partial_product_19(462) <= '0';
partial_product_19(463) <= '0';
partial_product_19(464) <= '0';
partial_product_19(465) <= '0';
partial_product_19(466) <= '0';
partial_product_19(467) <= '0';
partial_product_19(468) <= '0';
partial_product_19(469) <= '0';
partial_product_19(470) <= '0';
partial_product_19(471) <= '0';
partial_product_19(472) <= '0';
partial_product_19(473) <= '0';
partial_product_19(474) <= '0';
partial_product_19(475) <= '0';
partial_product_19(476) <= '0';
partial_product_19(477) <= '0';
partial_product_19(478) <= '0';
partial_product_19(479) <= '0';
partial_product_19(480) <= '0';
partial_product_19(481) <= '0';
partial_product_19(482) <= '0';
partial_product_19(483) <= '0';
partial_product_19(484) <= '0';
partial_product_19(485) <= '0';
partial_product_19(486) <= '0';
partial_product_19(487) <= '0';
partial_product_19(488) <= '0';
partial_product_19(489) <= '0';
partial_product_19(490) <= '0';
partial_product_19(491) <= '0';
partial_product_19(492) <= '0';
partial_product_19(493) <= '0';
partial_product_19(494) <= '0';
partial_product_19(495) <= '0';
partial_product_19(496) <= '0';
partial_product_19(497) <= '0';
partial_product_19(498) <= '0';
partial_product_19(499) <= '0';
partial_product_19(500) <= '0';
partial_product_19(501) <= '0';
partial_product_19(502) <= '0';
partial_product_19(503) <= '0';
partial_product_19(504) <= '0';
partial_product_19(505) <= '0';
partial_product_19(506) <= '0';
partial_product_19(507) <= '0';
partial_product_19(508) <= '0';
partial_product_19(509) <= '0';
partial_product_19(510) <= '0';
partial_product_19(511) <= '0';
partial_product_19(512) <= '0';
partial_product_20(0) <= '0';
partial_product_20(1) <= '0';
partial_product_20(2) <= '0';
partial_product_20(3) <= '0';
partial_product_20(4) <= '0';
partial_product_20(5) <= '0';
partial_product_20(6) <= '0';
partial_product_20(7) <= '0';
partial_product_20(8) <= '0';
partial_product_20(9) <= '0';
partial_product_20(10) <= '0';
partial_product_20(11) <= '0';
partial_product_20(12) <= '0';
partial_product_20(13) <= '0';
partial_product_20(14) <= '0';
partial_product_20(15) <= '0';
partial_product_20(16) <= '0';
partial_product_20(17) <= '0';
partial_product_20(18) <= '0';
partial_product_20(19) <= '0';
partial_product_20(20) <= '0';
partial_product_20(21) <= '0';
partial_product_20(22) <= '0';
partial_product_20(23) <= '0';
partial_product_20(24) <= '0';
partial_product_20(25) <= '0';
partial_product_20(26) <= '0';
partial_product_20(27) <= '0';
partial_product_20(28) <= '0';
partial_product_20(29) <= '0';
partial_product_20(30) <= '0';
partial_product_20(31) <= '0';
partial_product_20(32) <= '0';
partial_product_20(33) <= '0';
partial_product_20(34) <= '0';
partial_product_20(35) <= '0';
partial_product_20(36) <= '0';
partial_product_20(37) <= '0';
partial_product_20(38) <= '0';
partial_product_20(39) <= '0';
partial_product_20(40) <= '0';
partial_product_20(41) <= '0';
partial_product_20(42) <= '0';
partial_product_20(43) <= '0';
partial_product_20(44) <= '0';
partial_product_20(45) <= '0';
partial_product_20(46) <= '0';
partial_product_20(47) <= '0';
partial_product_20(48) <= '0';
partial_product_20(49) <= '0';
partial_product_20(50) <= '0';
partial_product_20(51) <= '0';
partial_product_20(52) <= '0';
partial_product_20(53) <= '0';
partial_product_20(54) <= '0';
partial_product_20(55) <= '0';
partial_product_20(56) <= '0';
partial_product_20(57) <= '0';
partial_product_20(58) <= '0';
partial_product_20(59) <= '0';
partial_product_20(60) <= '0';
partial_product_20(61) <= '0';
partial_product_20(62) <= '0';
partial_product_20(63) <= '0';
partial_product_20(64) <= '0';
partial_product_20(65) <= '0';
partial_product_20(66) <= '0';
partial_product_20(67) <= '0';
partial_product_20(68) <= '0';
partial_product_20(69) <= '0';
partial_product_20(70) <= '0';
partial_product_20(71) <= '0';
partial_product_20(72) <= '0';
partial_product_20(73) <= '0';
partial_product_20(74) <= '0';
partial_product_20(75) <= '0';
partial_product_20(76) <= '0';
partial_product_20(77) <= '0';
partial_product_20(78) <= '0';
partial_product_20(79) <= '0';
partial_product_20(80) <= '0';
partial_product_20(81) <= '0';
partial_product_20(82) <= '0';
partial_product_20(83) <= '0';
partial_product_20(84) <= '0';
partial_product_20(85) <= '0';
partial_product_20(86) <= '0';
partial_product_20(87) <= '0';
partial_product_20(88) <= '0';
partial_product_20(89) <= '0';
partial_product_20(90) <= '0';
partial_product_20(91) <= '0';
partial_product_20(92) <= '0';
partial_product_20(93) <= '0';
partial_product_20(94) <= '0';
partial_product_20(95) <= '0';
partial_product_20(96) <= '0';
partial_product_20(97) <= '0';
partial_product_20(98) <= '0';
partial_product_20(99) <= '0';
partial_product_20(100) <= '0';
partial_product_20(101) <= '0';
partial_product_20(102) <= '0';
partial_product_20(103) <= '0';
partial_product_20(104) <= '0';
partial_product_20(105) <= '0';
partial_product_20(106) <= '0';
partial_product_20(107) <= '0';
partial_product_20(108) <= '0';
partial_product_20(109) <= '0';
partial_product_20(110) <= '0';
partial_product_20(111) <= '0';
partial_product_20(112) <= '0';
partial_product_20(113) <= '0';
partial_product_20(114) <= '0';
partial_product_20(115) <= '0';
partial_product_20(116) <= '0';
partial_product_20(117) <= '0';
partial_product_20(118) <= '0';
partial_product_20(119) <= '0';
partial_product_20(120) <= '0';
partial_product_20(121) <= '0';
partial_product_20(122) <= '0';
partial_product_20(123) <= '0';
partial_product_20(124) <= '0';
partial_product_20(125) <= '0';
partial_product_20(126) <= '0';
partial_product_20(127) <= '0';
partial_product_20(128) <= '0';
partial_product_20(129) <= '0';
partial_product_20(130) <= '0';
partial_product_20(131) <= '0';
partial_product_20(132) <= '0';
partial_product_20(133) <= '0';
partial_product_20(134) <= '0';
partial_product_20(135) <= '0';
partial_product_20(136) <= '0';
partial_product_20(137) <= '0';
partial_product_20(138) <= '0';
partial_product_20(139) <= '0';
partial_product_20(140) <= '0';
partial_product_20(141) <= '0';
partial_product_20(142) <= '0';
partial_product_20(143) <= '0';
partial_product_20(144) <= '0';
partial_product_20(145) <= '0';
partial_product_20(146) <= '0';
partial_product_20(147) <= '0';
partial_product_20(148) <= '0';
partial_product_20(149) <= '0';
partial_product_20(150) <= '0';
partial_product_20(151) <= '0';
partial_product_20(152) <= '0';
partial_product_20(153) <= '0';
partial_product_20(154) <= '0';
partial_product_20(155) <= '0';
partial_product_20(156) <= '0';
partial_product_20(157) <= '0';
partial_product_20(158) <= '0';
partial_product_20(159) <= '0';
partial_product_20(160) <= '0';
partial_product_20(161) <= '0';
partial_product_20(162) <= '0';
partial_product_20(163) <= '0';
partial_product_20(164) <= '0';
partial_product_20(165) <= '0';
partial_product_20(166) <= '0';
partial_product_20(167) <= '0';
partial_product_20(168) <= '0';
partial_product_20(169) <= '0';
partial_product_20(170) <= '0';
partial_product_20(171) <= '0';
partial_product_20(172) <= '0';
partial_product_20(173) <= '0';
partial_product_20(174) <= '0';
partial_product_20(175) <= '0';
partial_product_20(176) <= '0';
partial_product_20(177) <= '0';
partial_product_20(178) <= '0';
partial_product_20(179) <= '0';
partial_product_20(180) <= '0';
partial_product_20(181) <= '0';
partial_product_20(182) <= '0';
partial_product_20(183) <= '0';
partial_product_20(184) <= '0';
partial_product_20(185) <= '0';
partial_product_20(186) <= '0';
partial_product_20(187) <= '0';
partial_product_20(188) <= '0';
partial_product_20(189) <= '0';
partial_product_20(190) <= '0';
partial_product_20(191) <= '0';
partial_product_20(192) <= '0';
partial_product_20(193) <= '0';
partial_product_20(194) <= '0';
partial_product_20(195) <= '0';
partial_product_20(196) <= '0';
partial_product_20(197) <= '0';
partial_product_20(198) <= '0';
partial_product_20(199) <= '0';
partial_product_20(200) <= '0';
partial_product_20(201) <= '0';
partial_product_20(202) <= '0';
partial_product_20(203) <= '0';
partial_product_20(204) <= temp_mult_84(204);
partial_product_20(205) <= temp_mult_84(205);
partial_product_20(206) <= temp_mult_84(206);
partial_product_20(207) <= temp_mult_84(207);
partial_product_20(208) <= temp_mult_84(208);
partial_product_20(209) <= temp_mult_84(209);
partial_product_20(210) <= temp_mult_84(210);
partial_product_20(211) <= temp_mult_84(211);
partial_product_20(212) <= temp_mult_84(212);
partial_product_20(213) <= temp_mult_84(213);
partial_product_20(214) <= temp_mult_84(214);
partial_product_20(215) <= temp_mult_84(215);
partial_product_20(216) <= temp_mult_84(216);
partial_product_20(217) <= temp_mult_84(217);
partial_product_20(218) <= temp_mult_84(218);
partial_product_20(219) <= temp_mult_84(219);
partial_product_20(220) <= temp_mult_84(220);
partial_product_20(221) <= temp_mult_84(221);
partial_product_20(222) <= temp_mult_84(222);
partial_product_20(223) <= temp_mult_84(223);
partial_product_20(224) <= temp_mult_84(224);
partial_product_20(225) <= temp_mult_84(225);
partial_product_20(226) <= temp_mult_84(226);
partial_product_20(227) <= temp_mult_84(227);
partial_product_20(228) <= temp_mult_84(228);
partial_product_20(229) <= temp_mult_84(229);
partial_product_20(230) <= temp_mult_84(230);
partial_product_20(231) <= temp_mult_84(231);
partial_product_20(232) <= temp_mult_84(232);
partial_product_20(233) <= temp_mult_84(233);
partial_product_20(234) <= temp_mult_84(234);
partial_product_20(235) <= temp_mult_84(235);
partial_product_20(236) <= temp_mult_84(236);
partial_product_20(237) <= temp_mult_84(237);
partial_product_20(238) <= temp_mult_84(238);
partial_product_20(239) <= temp_mult_84(239);
partial_product_20(240) <= temp_mult_84(240);
partial_product_20(241) <= temp_mult_84(241);
partial_product_20(242) <= temp_mult_84(242);
partial_product_20(243) <= temp_mult_84(243);
partial_product_20(244) <= temp_mult_84(244);
partial_product_20(245) <= temp_mult_93(245);
partial_product_20(246) <= temp_mult_93(246);
partial_product_20(247) <= temp_mult_93(247);
partial_product_20(248) <= temp_mult_93(248);
partial_product_20(249) <= temp_mult_93(249);
partial_product_20(250) <= temp_mult_93(250);
partial_product_20(251) <= temp_mult_93(251);
partial_product_20(252) <= temp_mult_93(252);
partial_product_20(253) <= temp_mult_93(253);
partial_product_20(254) <= temp_mult_93(254);
partial_product_20(255) <= temp_mult_93(255);
partial_product_20(256) <= temp_mult_93(256);
partial_product_20(257) <= temp_mult_93(257);
partial_product_20(258) <= temp_mult_93(258);
partial_product_20(259) <= temp_mult_93(259);
partial_product_20(260) <= temp_mult_93(260);
partial_product_20(261) <= temp_mult_93(261);
partial_product_20(262) <= temp_mult_93(262);
partial_product_20(263) <= temp_mult_93(263);
partial_product_20(264) <= temp_mult_93(264);
partial_product_20(265) <= temp_mult_93(265);
partial_product_20(266) <= temp_mult_93(266);
partial_product_20(267) <= temp_mult_93(267);
partial_product_20(268) <= temp_mult_93(268);
partial_product_20(269) <= temp_mult_93(269);
partial_product_20(270) <= temp_mult_93(270);
partial_product_20(271) <= temp_mult_93(271);
partial_product_20(272) <= temp_mult_93(272);
partial_product_20(273) <= temp_mult_93(273);
partial_product_20(274) <= temp_mult_93(274);
partial_product_20(275) <= temp_mult_93(275);
partial_product_20(276) <= temp_mult_93(276);
partial_product_20(277) <= temp_mult_93(277);
partial_product_20(278) <= temp_mult_93(278);
partial_product_20(279) <= temp_mult_93(279);
partial_product_20(280) <= temp_mult_93(280);
partial_product_20(281) <= temp_mult_93(281);
partial_product_20(282) <= temp_mult_93(282);
partial_product_20(283) <= temp_mult_93(283);
partial_product_20(284) <= temp_mult_93(284);
partial_product_20(285) <= temp_mult_93(285);
partial_product_20(286) <= temp_mult_102(286);
partial_product_20(287) <= temp_mult_102(287);
partial_product_20(288) <= temp_mult_102(288);
partial_product_20(289) <= temp_mult_102(289);
partial_product_20(290) <= temp_mult_102(290);
partial_product_20(291) <= temp_mult_102(291);
partial_product_20(292) <= temp_mult_102(292);
partial_product_20(293) <= temp_mult_102(293);
partial_product_20(294) <= temp_mult_102(294);
partial_product_20(295) <= temp_mult_102(295);
partial_product_20(296) <= temp_mult_102(296);
partial_product_20(297) <= temp_mult_102(297);
partial_product_20(298) <= temp_mult_102(298);
partial_product_20(299) <= temp_mult_102(299);
partial_product_20(300) <= temp_mult_102(300);
partial_product_20(301) <= temp_mult_102(301);
partial_product_20(302) <= temp_mult_102(302);
partial_product_20(303) <= temp_mult_102(303);
partial_product_20(304) <= temp_mult_102(304);
partial_product_20(305) <= temp_mult_102(305);
partial_product_20(306) <= temp_mult_102(306);
partial_product_20(307) <= temp_mult_102(307);
partial_product_20(308) <= temp_mult_102(308);
partial_product_20(309) <= temp_mult_102(309);
partial_product_20(310) <= temp_mult_102(310);
partial_product_20(311) <= temp_mult_102(311);
partial_product_20(312) <= temp_mult_102(312);
partial_product_20(313) <= temp_mult_102(313);
partial_product_20(314) <= temp_mult_102(314);
partial_product_20(315) <= temp_mult_102(315);
partial_product_20(316) <= temp_mult_102(316);
partial_product_20(317) <= temp_mult_102(317);
partial_product_20(318) <= temp_mult_102(318);
partial_product_20(319) <= temp_mult_102(319);
partial_product_20(320) <= temp_mult_102(320);
partial_product_20(321) <= temp_mult_102(321);
partial_product_20(322) <= temp_mult_102(322);
partial_product_20(323) <= temp_mult_102(323);
partial_product_20(324) <= temp_mult_102(324);
partial_product_20(325) <= temp_mult_102(325);
partial_product_20(326) <= temp_mult_102(326);
partial_product_20(327) <= '0';
partial_product_20(328) <= '0';
partial_product_20(329) <= '0';
partial_product_20(330) <= '0';
partial_product_20(331) <= '0';
partial_product_20(332) <= '0';
partial_product_20(333) <= '0';
partial_product_20(334) <= '0';
partial_product_20(335) <= '0';
partial_product_20(336) <= '0';
partial_product_20(337) <= '0';
partial_product_20(338) <= '0';
partial_product_20(339) <= '0';
partial_product_20(340) <= '0';
partial_product_20(341) <= '0';
partial_product_20(342) <= '0';
partial_product_20(343) <= '0';
partial_product_20(344) <= '0';
partial_product_20(345) <= '0';
partial_product_20(346) <= '0';
partial_product_20(347) <= '0';
partial_product_20(348) <= '0';
partial_product_20(349) <= '0';
partial_product_20(350) <= '0';
partial_product_20(351) <= '0';
partial_product_20(352) <= '0';
partial_product_20(353) <= '0';
partial_product_20(354) <= '0';
partial_product_20(355) <= '0';
partial_product_20(356) <= '0';
partial_product_20(357) <= '0';
partial_product_20(358) <= '0';
partial_product_20(359) <= '0';
partial_product_20(360) <= '0';
partial_product_20(361) <= '0';
partial_product_20(362) <= '0';
partial_product_20(363) <= '0';
partial_product_20(364) <= '0';
partial_product_20(365) <= '0';
partial_product_20(366) <= '0';
partial_product_20(367) <= '0';
partial_product_20(368) <= '0';
partial_product_20(369) <= '0';
partial_product_20(370) <= '0';
partial_product_20(371) <= '0';
partial_product_20(372) <= '0';
partial_product_20(373) <= '0';
partial_product_20(374) <= '0';
partial_product_20(375) <= '0';
partial_product_20(376) <= '0';
partial_product_20(377) <= '0';
partial_product_20(378) <= '0';
partial_product_20(379) <= '0';
partial_product_20(380) <= '0';
partial_product_20(381) <= '0';
partial_product_20(382) <= '0';
partial_product_20(383) <= '0';
partial_product_20(384) <= '0';
partial_product_20(385) <= '0';
partial_product_20(386) <= '0';
partial_product_20(387) <= '0';
partial_product_20(388) <= '0';
partial_product_20(389) <= '0';
partial_product_20(390) <= '0';
partial_product_20(391) <= '0';
partial_product_20(392) <= '0';
partial_product_20(393) <= '0';
partial_product_20(394) <= '0';
partial_product_20(395) <= '0';
partial_product_20(396) <= '0';
partial_product_20(397) <= '0';
partial_product_20(398) <= '0';
partial_product_20(399) <= '0';
partial_product_20(400) <= '0';
partial_product_20(401) <= '0';
partial_product_20(402) <= '0';
partial_product_20(403) <= '0';
partial_product_20(404) <= '0';
partial_product_20(405) <= '0';
partial_product_20(406) <= '0';
partial_product_20(407) <= '0';
partial_product_20(408) <= '0';
partial_product_20(409) <= '0';
partial_product_20(410) <= '0';
partial_product_20(411) <= '0';
partial_product_20(412) <= '0';
partial_product_20(413) <= '0';
partial_product_20(414) <= '0';
partial_product_20(415) <= '0';
partial_product_20(416) <= '0';
partial_product_20(417) <= '0';
partial_product_20(418) <= '0';
partial_product_20(419) <= '0';
partial_product_20(420) <= '0';
partial_product_20(421) <= '0';
partial_product_20(422) <= '0';
partial_product_20(423) <= '0';
partial_product_20(424) <= '0';
partial_product_20(425) <= '0';
partial_product_20(426) <= '0';
partial_product_20(427) <= '0';
partial_product_20(428) <= '0';
partial_product_20(429) <= '0';
partial_product_20(430) <= '0';
partial_product_20(431) <= '0';
partial_product_20(432) <= '0';
partial_product_20(433) <= '0';
partial_product_20(434) <= '0';
partial_product_20(435) <= '0';
partial_product_20(436) <= '0';
partial_product_20(437) <= '0';
partial_product_20(438) <= '0';
partial_product_20(439) <= '0';
partial_product_20(440) <= '0';
partial_product_20(441) <= '0';
partial_product_20(442) <= '0';
partial_product_20(443) <= '0';
partial_product_20(444) <= '0';
partial_product_20(445) <= '0';
partial_product_20(446) <= '0';
partial_product_20(447) <= '0';
partial_product_20(448) <= '0';
partial_product_20(449) <= '0';
partial_product_20(450) <= '0';
partial_product_20(451) <= '0';
partial_product_20(452) <= '0';
partial_product_20(453) <= '0';
partial_product_20(454) <= '0';
partial_product_20(455) <= '0';
partial_product_20(456) <= '0';
partial_product_20(457) <= '0';
partial_product_20(458) <= '0';
partial_product_20(459) <= '0';
partial_product_20(460) <= '0';
partial_product_20(461) <= '0';
partial_product_20(462) <= '0';
partial_product_20(463) <= '0';
partial_product_20(464) <= '0';
partial_product_20(465) <= '0';
partial_product_20(466) <= '0';
partial_product_20(467) <= '0';
partial_product_20(468) <= '0';
partial_product_20(469) <= '0';
partial_product_20(470) <= '0';
partial_product_20(471) <= '0';
partial_product_20(472) <= '0';
partial_product_20(473) <= '0';
partial_product_20(474) <= '0';
partial_product_20(475) <= '0';
partial_product_20(476) <= '0';
partial_product_20(477) <= '0';
partial_product_20(478) <= '0';
partial_product_20(479) <= '0';
partial_product_20(480) <= '0';
partial_product_20(481) <= '0';
partial_product_20(482) <= '0';
partial_product_20(483) <= '0';
partial_product_20(484) <= '0';
partial_product_20(485) <= '0';
partial_product_20(486) <= '0';
partial_product_20(487) <= '0';
partial_product_20(488) <= '0';
partial_product_20(489) <= '0';
partial_product_20(490) <= '0';
partial_product_20(491) <= '0';
partial_product_20(492) <= '0';
partial_product_20(493) <= '0';
partial_product_20(494) <= '0';
partial_product_20(495) <= '0';
partial_product_20(496) <= '0';
partial_product_20(497) <= '0';
partial_product_20(498) <= '0';
partial_product_20(499) <= '0';
partial_product_20(500) <= '0';
partial_product_20(501) <= '0';
partial_product_20(502) <= '0';
partial_product_20(503) <= '0';
partial_product_20(504) <= '0';
partial_product_20(505) <= '0';
partial_product_20(506) <= '0';
partial_product_20(507) <= '0';
partial_product_20(508) <= '0';
partial_product_20(509) <= '0';
partial_product_20(510) <= '0';
partial_product_20(511) <= '0';
partial_product_20(512) <= '0';
partial_product_21(0) <= '0';
partial_product_21(1) <= '0';
partial_product_21(2) <= '0';
partial_product_21(3) <= '0';
partial_product_21(4) <= '0';
partial_product_21(5) <= '0';
partial_product_21(6) <= '0';
partial_product_21(7) <= '0';
partial_product_21(8) <= '0';
partial_product_21(9) <= '0';
partial_product_21(10) <= '0';
partial_product_21(11) <= '0';
partial_product_21(12) <= '0';
partial_product_21(13) <= '0';
partial_product_21(14) <= '0';
partial_product_21(15) <= '0';
partial_product_21(16) <= '0';
partial_product_21(17) <= '0';
partial_product_21(18) <= '0';
partial_product_21(19) <= '0';
partial_product_21(20) <= '0';
partial_product_21(21) <= '0';
partial_product_21(22) <= '0';
partial_product_21(23) <= '0';
partial_product_21(24) <= '0';
partial_product_21(25) <= '0';
partial_product_21(26) <= '0';
partial_product_21(27) <= '0';
partial_product_21(28) <= '0';
partial_product_21(29) <= '0';
partial_product_21(30) <= '0';
partial_product_21(31) <= '0';
partial_product_21(32) <= '0';
partial_product_21(33) <= '0';
partial_product_21(34) <= '0';
partial_product_21(35) <= '0';
partial_product_21(36) <= '0';
partial_product_21(37) <= '0';
partial_product_21(38) <= '0';
partial_product_21(39) <= '0';
partial_product_21(40) <= '0';
partial_product_21(41) <= '0';
partial_product_21(42) <= '0';
partial_product_21(43) <= '0';
partial_product_21(44) <= '0';
partial_product_21(45) <= '0';
partial_product_21(46) <= '0';
partial_product_21(47) <= '0';
partial_product_21(48) <= '0';
partial_product_21(49) <= '0';
partial_product_21(50) <= '0';
partial_product_21(51) <= '0';
partial_product_21(52) <= '0';
partial_product_21(53) <= '0';
partial_product_21(54) <= '0';
partial_product_21(55) <= '0';
partial_product_21(56) <= '0';
partial_product_21(57) <= '0';
partial_product_21(58) <= '0';
partial_product_21(59) <= '0';
partial_product_21(60) <= '0';
partial_product_21(61) <= '0';
partial_product_21(62) <= '0';
partial_product_21(63) <= '0';
partial_product_21(64) <= '0';
partial_product_21(65) <= '0';
partial_product_21(66) <= '0';
partial_product_21(67) <= '0';
partial_product_21(68) <= '0';
partial_product_21(69) <= '0';
partial_product_21(70) <= '0';
partial_product_21(71) <= '0';
partial_product_21(72) <= '0';
partial_product_21(73) <= '0';
partial_product_21(74) <= '0';
partial_product_21(75) <= '0';
partial_product_21(76) <= '0';
partial_product_21(77) <= '0';
partial_product_21(78) <= '0';
partial_product_21(79) <= '0';
partial_product_21(80) <= '0';
partial_product_21(81) <= '0';
partial_product_21(82) <= '0';
partial_product_21(83) <= '0';
partial_product_21(84) <= '0';
partial_product_21(85) <= '0';
partial_product_21(86) <= '0';
partial_product_21(87) <= '0';
partial_product_21(88) <= '0';
partial_product_21(89) <= '0';
partial_product_21(90) <= '0';
partial_product_21(91) <= '0';
partial_product_21(92) <= '0';
partial_product_21(93) <= '0';
partial_product_21(94) <= '0';
partial_product_21(95) <= '0';
partial_product_21(96) <= '0';
partial_product_21(97) <= '0';
partial_product_21(98) <= '0';
partial_product_21(99) <= '0';
partial_product_21(100) <= '0';
partial_product_21(101) <= '0';
partial_product_21(102) <= '0';
partial_product_21(103) <= '0';
partial_product_21(104) <= '0';
partial_product_21(105) <= '0';
partial_product_21(106) <= '0';
partial_product_21(107) <= '0';
partial_product_21(108) <= '0';
partial_product_21(109) <= '0';
partial_product_21(110) <= '0';
partial_product_21(111) <= '0';
partial_product_21(112) <= '0';
partial_product_21(113) <= '0';
partial_product_21(114) <= '0';
partial_product_21(115) <= '0';
partial_product_21(116) <= '0';
partial_product_21(117) <= '0';
partial_product_21(118) <= '0';
partial_product_21(119) <= '0';
partial_product_21(120) <= '0';
partial_product_21(121) <= '0';
partial_product_21(122) <= '0';
partial_product_21(123) <= '0';
partial_product_21(124) <= '0';
partial_product_21(125) <= '0';
partial_product_21(126) <= '0';
partial_product_21(127) <= '0';
partial_product_21(128) <= '0';
partial_product_21(129) <= '0';
partial_product_21(130) <= '0';
partial_product_21(131) <= '0';
partial_product_21(132) <= '0';
partial_product_21(133) <= '0';
partial_product_21(134) <= '0';
partial_product_21(135) <= '0';
partial_product_21(136) <= '0';
partial_product_21(137) <= '0';
partial_product_21(138) <= '0';
partial_product_21(139) <= '0';
partial_product_21(140) <= '0';
partial_product_21(141) <= '0';
partial_product_21(142) <= '0';
partial_product_21(143) <= '0';
partial_product_21(144) <= '0';
partial_product_21(145) <= '0';
partial_product_21(146) <= '0';
partial_product_21(147) <= '0';
partial_product_21(148) <= '0';
partial_product_21(149) <= '0';
partial_product_21(150) <= '0';
partial_product_21(151) <= '0';
partial_product_21(152) <= '0';
partial_product_21(153) <= '0';
partial_product_21(154) <= '0';
partial_product_21(155) <= '0';
partial_product_21(156) <= '0';
partial_product_21(157) <= '0';
partial_product_21(158) <= '0';
partial_product_21(159) <= '0';
partial_product_21(160) <= '0';
partial_product_21(161) <= '0';
partial_product_21(162) <= '0';
partial_product_21(163) <= '0';
partial_product_21(164) <= '0';
partial_product_21(165) <= '0';
partial_product_21(166) <= '0';
partial_product_21(167) <= '0';
partial_product_21(168) <= '0';
partial_product_21(169) <= '0';
partial_product_21(170) <= '0';
partial_product_21(171) <= '0';
partial_product_21(172) <= '0';
partial_product_21(173) <= '0';
partial_product_21(174) <= '0';
partial_product_21(175) <= '0';
partial_product_21(176) <= '0';
partial_product_21(177) <= '0';
partial_product_21(178) <= '0';
partial_product_21(179) <= '0';
partial_product_21(180) <= '0';
partial_product_21(181) <= '0';
partial_product_21(182) <= '0';
partial_product_21(183) <= '0';
partial_product_21(184) <= '0';
partial_product_21(185) <= '0';
partial_product_21(186) <= '0';
partial_product_21(187) <= '0';
partial_product_21(188) <= '0';
partial_product_21(189) <= '0';
partial_product_21(190) <= '0';
partial_product_21(191) <= '0';
partial_product_21(192) <= '0';
partial_product_21(193) <= '0';
partial_product_21(194) <= '0';
partial_product_21(195) <= '0';
partial_product_21(196) <= '0';
partial_product_21(197) <= '0';
partial_product_21(198) <= '0';
partial_product_21(199) <= '0';
partial_product_21(200) <= '0';
partial_product_21(201) <= '0';
partial_product_21(202) <= '0';
partial_product_21(203) <= '0';
partial_product_21(204) <= '0';
partial_product_21(205) <= '0';
partial_product_21(206) <= '0';
partial_product_21(207) <= '0';
partial_product_21(208) <= '0';
partial_product_21(209) <= '0';
partial_product_21(210) <= '0';
partial_product_21(211) <= '0';
partial_product_21(212) <= '0';
partial_product_21(213) <= '0';
partial_product_21(214) <= '0';
partial_product_21(215) <= '0';
partial_product_21(216) <= temp_mult_72(216);
partial_product_21(217) <= temp_mult_72(217);
partial_product_21(218) <= temp_mult_72(218);
partial_product_21(219) <= temp_mult_72(219);
partial_product_21(220) <= temp_mult_72(220);
partial_product_21(221) <= temp_mult_72(221);
partial_product_21(222) <= temp_mult_72(222);
partial_product_21(223) <= temp_mult_72(223);
partial_product_21(224) <= temp_mult_72(224);
partial_product_21(225) <= temp_mult_72(225);
partial_product_21(226) <= temp_mult_72(226);
partial_product_21(227) <= temp_mult_72(227);
partial_product_21(228) <= temp_mult_72(228);
partial_product_21(229) <= temp_mult_72(229);
partial_product_21(230) <= temp_mult_72(230);
partial_product_21(231) <= temp_mult_72(231);
partial_product_21(232) <= temp_mult_72(232);
partial_product_21(233) <= temp_mult_72(233);
partial_product_21(234) <= temp_mult_72(234);
partial_product_21(235) <= temp_mult_72(235);
partial_product_21(236) <= temp_mult_72(236);
partial_product_21(237) <= temp_mult_72(237);
partial_product_21(238) <= temp_mult_72(238);
partial_product_21(239) <= temp_mult_72(239);
partial_product_21(240) <= temp_mult_72(240);
partial_product_21(241) <= temp_mult_72(241);
partial_product_21(242) <= temp_mult_72(242);
partial_product_21(243) <= temp_mult_72(243);
partial_product_21(244) <= temp_mult_72(244);
partial_product_21(245) <= temp_mult_72(245);
partial_product_21(246) <= temp_mult_72(246);
partial_product_21(247) <= temp_mult_72(247);
partial_product_21(248) <= temp_mult_72(248);
partial_product_21(249) <= temp_mult_72(249);
partial_product_21(250) <= temp_mult_72(250);
partial_product_21(251) <= temp_mult_72(251);
partial_product_21(252) <= temp_mult_72(252);
partial_product_21(253) <= temp_mult_72(253);
partial_product_21(254) <= temp_mult_72(254);
partial_product_21(255) <= temp_mult_72(255);
partial_product_21(256) <= temp_mult_72(256);
partial_product_21(257) <= '0';
partial_product_21(258) <= '0';
partial_product_21(259) <= '0';
partial_product_21(260) <= '0';
partial_product_21(261) <= '0';
partial_product_21(262) <= temp_mult_94(262);
partial_product_21(263) <= temp_mult_94(263);
partial_product_21(264) <= temp_mult_94(264);
partial_product_21(265) <= temp_mult_94(265);
partial_product_21(266) <= temp_mult_94(266);
partial_product_21(267) <= temp_mult_94(267);
partial_product_21(268) <= temp_mult_94(268);
partial_product_21(269) <= temp_mult_94(269);
partial_product_21(270) <= temp_mult_94(270);
partial_product_21(271) <= temp_mult_94(271);
partial_product_21(272) <= temp_mult_94(272);
partial_product_21(273) <= temp_mult_94(273);
partial_product_21(274) <= temp_mult_94(274);
partial_product_21(275) <= temp_mult_94(275);
partial_product_21(276) <= temp_mult_94(276);
partial_product_21(277) <= temp_mult_94(277);
partial_product_21(278) <= temp_mult_94(278);
partial_product_21(279) <= temp_mult_94(279);
partial_product_21(280) <= temp_mult_94(280);
partial_product_21(281) <= temp_mult_94(281);
partial_product_21(282) <= temp_mult_94(282);
partial_product_21(283) <= temp_mult_94(283);
partial_product_21(284) <= temp_mult_94(284);
partial_product_21(285) <= temp_mult_94(285);
partial_product_21(286) <= temp_mult_94(286);
partial_product_21(287) <= temp_mult_94(287);
partial_product_21(288) <= temp_mult_94(288);
partial_product_21(289) <= temp_mult_94(289);
partial_product_21(290) <= temp_mult_94(290);
partial_product_21(291) <= temp_mult_94(291);
partial_product_21(292) <= temp_mult_94(292);
partial_product_21(293) <= temp_mult_94(293);
partial_product_21(294) <= temp_mult_94(294);
partial_product_21(295) <= temp_mult_94(295);
partial_product_21(296) <= temp_mult_94(296);
partial_product_21(297) <= temp_mult_94(297);
partial_product_21(298) <= temp_mult_94(298);
partial_product_21(299) <= temp_mult_94(299);
partial_product_21(300) <= temp_mult_94(300);
partial_product_21(301) <= temp_mult_94(301);
partial_product_21(302) <= temp_mult_94(302);
partial_product_21(303) <= '0';
partial_product_21(304) <= '0';
partial_product_21(305) <= '0';
partial_product_21(306) <= '0';
partial_product_21(307) <= '0';
partial_product_21(308) <= '0';
partial_product_21(309) <= '0';
partial_product_21(310) <= '0';
partial_product_21(311) <= '0';
partial_product_21(312) <= '0';
partial_product_21(313) <= '0';
partial_product_21(314) <= '0';
partial_product_21(315) <= '0';
partial_product_21(316) <= '0';
partial_product_21(317) <= '0';
partial_product_21(318) <= '0';
partial_product_21(319) <= '0';
partial_product_21(320) <= '0';
partial_product_21(321) <= '0';
partial_product_21(322) <= '0';
partial_product_21(323) <= '0';
partial_product_21(324) <= '0';
partial_product_21(325) <= '0';
partial_product_21(326) <= '0';
partial_product_21(327) <= '0';
partial_product_21(328) <= '0';
partial_product_21(329) <= '0';
partial_product_21(330) <= '0';
partial_product_21(331) <= '0';
partial_product_21(332) <= '0';
partial_product_21(333) <= '0';
partial_product_21(334) <= '0';
partial_product_21(335) <= '0';
partial_product_21(336) <= '0';
partial_product_21(337) <= '0';
partial_product_21(338) <= '0';
partial_product_21(339) <= '0';
partial_product_21(340) <= '0';
partial_product_21(341) <= '0';
partial_product_21(342) <= '0';
partial_product_21(343) <= '0';
partial_product_21(344) <= '0';
partial_product_21(345) <= '0';
partial_product_21(346) <= '0';
partial_product_21(347) <= '0';
partial_product_21(348) <= '0';
partial_product_21(349) <= '0';
partial_product_21(350) <= '0';
partial_product_21(351) <= '0';
partial_product_21(352) <= '0';
partial_product_21(353) <= '0';
partial_product_21(354) <= '0';
partial_product_21(355) <= '0';
partial_product_21(356) <= '0';
partial_product_21(357) <= '0';
partial_product_21(358) <= '0';
partial_product_21(359) <= '0';
partial_product_21(360) <= '0';
partial_product_21(361) <= '0';
partial_product_21(362) <= '0';
partial_product_21(363) <= '0';
partial_product_21(364) <= '0';
partial_product_21(365) <= '0';
partial_product_21(366) <= '0';
partial_product_21(367) <= '0';
partial_product_21(368) <= '0';
partial_product_21(369) <= '0';
partial_product_21(370) <= '0';
partial_product_21(371) <= '0';
partial_product_21(372) <= '0';
partial_product_21(373) <= '0';
partial_product_21(374) <= '0';
partial_product_21(375) <= '0';
partial_product_21(376) <= '0';
partial_product_21(377) <= '0';
partial_product_21(378) <= '0';
partial_product_21(379) <= '0';
partial_product_21(380) <= '0';
partial_product_21(381) <= '0';
partial_product_21(382) <= '0';
partial_product_21(383) <= '0';
partial_product_21(384) <= '0';
partial_product_21(385) <= '0';
partial_product_21(386) <= '0';
partial_product_21(387) <= '0';
partial_product_21(388) <= '0';
partial_product_21(389) <= '0';
partial_product_21(390) <= '0';
partial_product_21(391) <= '0';
partial_product_21(392) <= '0';
partial_product_21(393) <= '0';
partial_product_21(394) <= '0';
partial_product_21(395) <= '0';
partial_product_21(396) <= '0';
partial_product_21(397) <= '0';
partial_product_21(398) <= '0';
partial_product_21(399) <= '0';
partial_product_21(400) <= '0';
partial_product_21(401) <= '0';
partial_product_21(402) <= '0';
partial_product_21(403) <= '0';
partial_product_21(404) <= '0';
partial_product_21(405) <= '0';
partial_product_21(406) <= '0';
partial_product_21(407) <= '0';
partial_product_21(408) <= '0';
partial_product_21(409) <= '0';
partial_product_21(410) <= '0';
partial_product_21(411) <= '0';
partial_product_21(412) <= '0';
partial_product_21(413) <= '0';
partial_product_21(414) <= '0';
partial_product_21(415) <= '0';
partial_product_21(416) <= '0';
partial_product_21(417) <= '0';
partial_product_21(418) <= '0';
partial_product_21(419) <= '0';
partial_product_21(420) <= '0';
partial_product_21(421) <= '0';
partial_product_21(422) <= '0';
partial_product_21(423) <= '0';
partial_product_21(424) <= '0';
partial_product_21(425) <= '0';
partial_product_21(426) <= '0';
partial_product_21(427) <= '0';
partial_product_21(428) <= '0';
partial_product_21(429) <= '0';
partial_product_21(430) <= '0';
partial_product_21(431) <= '0';
partial_product_21(432) <= '0';
partial_product_21(433) <= '0';
partial_product_21(434) <= '0';
partial_product_21(435) <= '0';
partial_product_21(436) <= '0';
partial_product_21(437) <= '0';
partial_product_21(438) <= '0';
partial_product_21(439) <= '0';
partial_product_21(440) <= '0';
partial_product_21(441) <= '0';
partial_product_21(442) <= '0';
partial_product_21(443) <= '0';
partial_product_21(444) <= '0';
partial_product_21(445) <= '0';
partial_product_21(446) <= '0';
partial_product_21(447) <= '0';
partial_product_21(448) <= '0';
partial_product_21(449) <= '0';
partial_product_21(450) <= '0';
partial_product_21(451) <= '0';
partial_product_21(452) <= '0';
partial_product_21(453) <= '0';
partial_product_21(454) <= '0';
partial_product_21(455) <= '0';
partial_product_21(456) <= '0';
partial_product_21(457) <= '0';
partial_product_21(458) <= '0';
partial_product_21(459) <= '0';
partial_product_21(460) <= '0';
partial_product_21(461) <= '0';
partial_product_21(462) <= '0';
partial_product_21(463) <= '0';
partial_product_21(464) <= '0';
partial_product_21(465) <= '0';
partial_product_21(466) <= '0';
partial_product_21(467) <= '0';
partial_product_21(468) <= '0';
partial_product_21(469) <= '0';
partial_product_21(470) <= '0';
partial_product_21(471) <= '0';
partial_product_21(472) <= '0';
partial_product_21(473) <= '0';
partial_product_21(474) <= '0';
partial_product_21(475) <= '0';
partial_product_21(476) <= '0';
partial_product_21(477) <= '0';
partial_product_21(478) <= '0';
partial_product_21(479) <= '0';
partial_product_21(480) <= '0';
partial_product_21(481) <= '0';
partial_product_21(482) <= '0';
partial_product_21(483) <= '0';
partial_product_21(484) <= '0';
partial_product_21(485) <= '0';
partial_product_21(486) <= '0';
partial_product_21(487) <= '0';
partial_product_21(488) <= '0';
partial_product_21(489) <= '0';
partial_product_21(490) <= '0';
partial_product_21(491) <= '0';
partial_product_21(492) <= '0';
partial_product_21(493) <= '0';
partial_product_21(494) <= '0';
partial_product_21(495) <= '0';
partial_product_21(496) <= '0';
partial_product_21(497) <= '0';
partial_product_21(498) <= '0';
partial_product_21(499) <= '0';
partial_product_21(500) <= '0';
partial_product_21(501) <= '0';
partial_product_21(502) <= '0';
partial_product_21(503) <= '0';
partial_product_21(504) <= '0';
partial_product_21(505) <= '0';
partial_product_21(506) <= '0';
partial_product_21(507) <= '0';
partial_product_21(508) <= '0';
partial_product_21(509) <= '0';
partial_product_21(510) <= '0';
partial_product_21(511) <= '0';
partial_product_21(512) <= '0';
partial_product_22(0) <= '0';
partial_product_22(1) <= '0';
partial_product_22(2) <= '0';
partial_product_22(3) <= '0';
partial_product_22(4) <= '0';
partial_product_22(5) <= '0';
partial_product_22(6) <= '0';
partial_product_22(7) <= '0';
partial_product_22(8) <= '0';
partial_product_22(9) <= '0';
partial_product_22(10) <= '0';
partial_product_22(11) <= '0';
partial_product_22(12) <= '0';
partial_product_22(13) <= '0';
partial_product_22(14) <= '0';
partial_product_22(15) <= '0';
partial_product_22(16) <= '0';
partial_product_22(17) <= '0';
partial_product_22(18) <= '0';
partial_product_22(19) <= '0';
partial_product_22(20) <= '0';
partial_product_22(21) <= '0';
partial_product_22(22) <= '0';
partial_product_22(23) <= '0';
partial_product_22(24) <= '0';
partial_product_22(25) <= '0';
partial_product_22(26) <= '0';
partial_product_22(27) <= '0';
partial_product_22(28) <= '0';
partial_product_22(29) <= '0';
partial_product_22(30) <= '0';
partial_product_22(31) <= '0';
partial_product_22(32) <= '0';
partial_product_22(33) <= '0';
partial_product_22(34) <= '0';
partial_product_22(35) <= '0';
partial_product_22(36) <= '0';
partial_product_22(37) <= '0';
partial_product_22(38) <= '0';
partial_product_22(39) <= '0';
partial_product_22(40) <= '0';
partial_product_22(41) <= '0';
partial_product_22(42) <= '0';
partial_product_22(43) <= '0';
partial_product_22(44) <= '0';
partial_product_22(45) <= '0';
partial_product_22(46) <= '0';
partial_product_22(47) <= '0';
partial_product_22(48) <= '0';
partial_product_22(49) <= '0';
partial_product_22(50) <= '0';
partial_product_22(51) <= '0';
partial_product_22(52) <= '0';
partial_product_22(53) <= '0';
partial_product_22(54) <= '0';
partial_product_22(55) <= '0';
partial_product_22(56) <= '0';
partial_product_22(57) <= '0';
partial_product_22(58) <= '0';
partial_product_22(59) <= '0';
partial_product_22(60) <= '0';
partial_product_22(61) <= '0';
partial_product_22(62) <= '0';
partial_product_22(63) <= '0';
partial_product_22(64) <= '0';
partial_product_22(65) <= '0';
partial_product_22(66) <= '0';
partial_product_22(67) <= '0';
partial_product_22(68) <= '0';
partial_product_22(69) <= '0';
partial_product_22(70) <= '0';
partial_product_22(71) <= '0';
partial_product_22(72) <= '0';
partial_product_22(73) <= '0';
partial_product_22(74) <= '0';
partial_product_22(75) <= '0';
partial_product_22(76) <= '0';
partial_product_22(77) <= '0';
partial_product_22(78) <= '0';
partial_product_22(79) <= '0';
partial_product_22(80) <= '0';
partial_product_22(81) <= '0';
partial_product_22(82) <= '0';
partial_product_22(83) <= '0';
partial_product_22(84) <= '0';
partial_product_22(85) <= '0';
partial_product_22(86) <= '0';
partial_product_22(87) <= '0';
partial_product_22(88) <= '0';
partial_product_22(89) <= '0';
partial_product_22(90) <= '0';
partial_product_22(91) <= '0';
partial_product_22(92) <= '0';
partial_product_22(93) <= '0';
partial_product_22(94) <= '0';
partial_product_22(95) <= '0';
partial_product_22(96) <= '0';
partial_product_22(97) <= '0';
partial_product_22(98) <= '0';
partial_product_22(99) <= '0';
partial_product_22(100) <= '0';
partial_product_22(101) <= '0';
partial_product_22(102) <= '0';
partial_product_22(103) <= '0';
partial_product_22(104) <= '0';
partial_product_22(105) <= '0';
partial_product_22(106) <= '0';
partial_product_22(107) <= '0';
partial_product_22(108) <= '0';
partial_product_22(109) <= '0';
partial_product_22(110) <= '0';
partial_product_22(111) <= '0';
partial_product_22(112) <= '0';
partial_product_22(113) <= '0';
partial_product_22(114) <= '0';
partial_product_22(115) <= '0';
partial_product_22(116) <= '0';
partial_product_22(117) <= '0';
partial_product_22(118) <= '0';
partial_product_22(119) <= '0';
partial_product_22(120) <= '0';
partial_product_22(121) <= '0';
partial_product_22(122) <= '0';
partial_product_22(123) <= '0';
partial_product_22(124) <= '0';
partial_product_22(125) <= '0';
partial_product_22(126) <= '0';
partial_product_22(127) <= '0';
partial_product_22(128) <= '0';
partial_product_22(129) <= '0';
partial_product_22(130) <= '0';
partial_product_22(131) <= '0';
partial_product_22(132) <= '0';
partial_product_22(133) <= '0';
partial_product_22(134) <= '0';
partial_product_22(135) <= '0';
partial_product_22(136) <= '0';
partial_product_22(137) <= '0';
partial_product_22(138) <= '0';
partial_product_22(139) <= '0';
partial_product_22(140) <= '0';
partial_product_22(141) <= '0';
partial_product_22(142) <= '0';
partial_product_22(143) <= '0';
partial_product_22(144) <= '0';
partial_product_22(145) <= '0';
partial_product_22(146) <= '0';
partial_product_22(147) <= '0';
partial_product_22(148) <= '0';
partial_product_22(149) <= '0';
partial_product_22(150) <= '0';
partial_product_22(151) <= '0';
partial_product_22(152) <= '0';
partial_product_22(153) <= '0';
partial_product_22(154) <= '0';
partial_product_22(155) <= '0';
partial_product_22(156) <= '0';
partial_product_22(157) <= '0';
partial_product_22(158) <= '0';
partial_product_22(159) <= '0';
partial_product_22(160) <= '0';
partial_product_22(161) <= '0';
partial_product_22(162) <= '0';
partial_product_22(163) <= '0';
partial_product_22(164) <= '0';
partial_product_22(165) <= '0';
partial_product_22(166) <= '0';
partial_product_22(167) <= '0';
partial_product_22(168) <= '0';
partial_product_22(169) <= '0';
partial_product_22(170) <= '0';
partial_product_22(171) <= '0';
partial_product_22(172) <= '0';
partial_product_22(173) <= '0';
partial_product_22(174) <= '0';
partial_product_22(175) <= '0';
partial_product_22(176) <= '0';
partial_product_22(177) <= '0';
partial_product_22(178) <= '0';
partial_product_22(179) <= '0';
partial_product_22(180) <= '0';
partial_product_22(181) <= '0';
partial_product_22(182) <= '0';
partial_product_22(183) <= '0';
partial_product_22(184) <= '0';
partial_product_22(185) <= '0';
partial_product_22(186) <= '0';
partial_product_22(187) <= '0';
partial_product_22(188) <= '0';
partial_product_22(189) <= '0';
partial_product_22(190) <= '0';
partial_product_22(191) <= '0';
partial_product_22(192) <= '0';
partial_product_22(193) <= '0';
partial_product_22(194) <= '0';
partial_product_22(195) <= '0';
partial_product_22(196) <= '0';
partial_product_22(197) <= '0';
partial_product_22(198) <= '0';
partial_product_22(199) <= '0';
partial_product_22(200) <= '0';
partial_product_22(201) <= '0';
partial_product_22(202) <= '0';
partial_product_22(203) <= '0';
partial_product_22(204) <= '0';
partial_product_22(205) <= '0';
partial_product_22(206) <= '0';
partial_product_22(207) <= '0';
partial_product_22(208) <= '0';
partial_product_22(209) <= '0';
partial_product_22(210) <= '0';
partial_product_22(211) <= '0';
partial_product_22(212) <= '0';
partial_product_22(213) <= '0';
partial_product_22(214) <= '0';
partial_product_22(215) <= '0';
partial_product_22(216) <= '0';
partial_product_22(217) <= '0';
partial_product_22(218) <= '0';
partial_product_22(219) <= '0';
partial_product_22(220) <= '0';
partial_product_22(221) <= temp_mult_85(221);
partial_product_22(222) <= temp_mult_85(222);
partial_product_22(223) <= temp_mult_85(223);
partial_product_22(224) <= temp_mult_85(224);
partial_product_22(225) <= temp_mult_85(225);
partial_product_22(226) <= temp_mult_85(226);
partial_product_22(227) <= temp_mult_85(227);
partial_product_22(228) <= temp_mult_85(228);
partial_product_22(229) <= temp_mult_85(229);
partial_product_22(230) <= temp_mult_85(230);
partial_product_22(231) <= temp_mult_85(231);
partial_product_22(232) <= temp_mult_85(232);
partial_product_22(233) <= temp_mult_85(233);
partial_product_22(234) <= temp_mult_85(234);
partial_product_22(235) <= temp_mult_85(235);
partial_product_22(236) <= temp_mult_85(236);
partial_product_22(237) <= temp_mult_85(237);
partial_product_22(238) <= temp_mult_85(238);
partial_product_22(239) <= temp_mult_85(239);
partial_product_22(240) <= temp_mult_85(240);
partial_product_22(241) <= temp_mult_85(241);
partial_product_22(242) <= temp_mult_85(242);
partial_product_22(243) <= temp_mult_85(243);
partial_product_22(244) <= temp_mult_85(244);
partial_product_22(245) <= temp_mult_85(245);
partial_product_22(246) <= temp_mult_85(246);
partial_product_22(247) <= temp_mult_85(247);
partial_product_22(248) <= temp_mult_85(248);
partial_product_22(249) <= temp_mult_85(249);
partial_product_22(250) <= temp_mult_85(250);
partial_product_22(251) <= temp_mult_85(251);
partial_product_22(252) <= temp_mult_85(252);
partial_product_22(253) <= temp_mult_85(253);
partial_product_22(254) <= temp_mult_85(254);
partial_product_22(255) <= temp_mult_85(255);
partial_product_22(256) <= temp_mult_85(256);
partial_product_22(257) <= temp_mult_85(257);
partial_product_22(258) <= temp_mult_85(258);
partial_product_22(259) <= temp_mult_85(259);
partial_product_22(260) <= temp_mult_85(260);
partial_product_22(261) <= temp_mult_85(261);
partial_product_22(262) <= '0';
partial_product_22(263) <= '0';
partial_product_22(264) <= '0';
partial_product_22(265) <= '0';
partial_product_22(266) <= '0';
partial_product_22(267) <= '0';
partial_product_22(268) <= '0';
partial_product_22(269) <= '0';
partial_product_22(270) <= '0';
partial_product_22(271) <= '0';
partial_product_22(272) <= '0';
partial_product_22(273) <= '0';
partial_product_22(274) <= '0';
partial_product_22(275) <= '0';
partial_product_22(276) <= '0';
partial_product_22(277) <= '0';
partial_product_22(278) <= '0';
partial_product_22(279) <= '0';
partial_product_22(280) <= '0';
partial_product_22(281) <= '0';
partial_product_22(282) <= '0';
partial_product_22(283) <= '0';
partial_product_22(284) <= '0';
partial_product_22(285) <= '0';
partial_product_22(286) <= '0';
partial_product_22(287) <= '0';
partial_product_22(288) <= '0';
partial_product_22(289) <= '0';
partial_product_22(290) <= '0';
partial_product_22(291) <= '0';
partial_product_22(292) <= '0';
partial_product_22(293) <= '0';
partial_product_22(294) <= '0';
partial_product_22(295) <= '0';
partial_product_22(296) <= '0';
partial_product_22(297) <= '0';
partial_product_22(298) <= '0';
partial_product_22(299) <= '0';
partial_product_22(300) <= '0';
partial_product_22(301) <= '0';
partial_product_22(302) <= '0';
partial_product_22(303) <= '0';
partial_product_22(304) <= '0';
partial_product_22(305) <= '0';
partial_product_22(306) <= '0';
partial_product_22(307) <= '0';
partial_product_22(308) <= '0';
partial_product_22(309) <= '0';
partial_product_22(310) <= '0';
partial_product_22(311) <= '0';
partial_product_22(312) <= '0';
partial_product_22(313) <= '0';
partial_product_22(314) <= '0';
partial_product_22(315) <= '0';
partial_product_22(316) <= '0';
partial_product_22(317) <= '0';
partial_product_22(318) <= '0';
partial_product_22(319) <= '0';
partial_product_22(320) <= '0';
partial_product_22(321) <= '0';
partial_product_22(322) <= '0';
partial_product_22(323) <= '0';
partial_product_22(324) <= '0';
partial_product_22(325) <= '0';
partial_product_22(326) <= '0';
partial_product_22(327) <= '0';
partial_product_22(328) <= '0';
partial_product_22(329) <= '0';
partial_product_22(330) <= '0';
partial_product_22(331) <= '0';
partial_product_22(332) <= '0';
partial_product_22(333) <= '0';
partial_product_22(334) <= '0';
partial_product_22(335) <= '0';
partial_product_22(336) <= '0';
partial_product_22(337) <= '0';
partial_product_22(338) <= '0';
partial_product_22(339) <= '0';
partial_product_22(340) <= '0';
partial_product_22(341) <= '0';
partial_product_22(342) <= '0';
partial_product_22(343) <= '0';
partial_product_22(344) <= '0';
partial_product_22(345) <= '0';
partial_product_22(346) <= '0';
partial_product_22(347) <= '0';
partial_product_22(348) <= '0';
partial_product_22(349) <= '0';
partial_product_22(350) <= '0';
partial_product_22(351) <= '0';
partial_product_22(352) <= '0';
partial_product_22(353) <= '0';
partial_product_22(354) <= '0';
partial_product_22(355) <= '0';
partial_product_22(356) <= '0';
partial_product_22(357) <= '0';
partial_product_22(358) <= '0';
partial_product_22(359) <= '0';
partial_product_22(360) <= '0';
partial_product_22(361) <= '0';
partial_product_22(362) <= '0';
partial_product_22(363) <= '0';
partial_product_22(364) <= '0';
partial_product_22(365) <= '0';
partial_product_22(366) <= '0';
partial_product_22(367) <= '0';
partial_product_22(368) <= '0';
partial_product_22(369) <= '0';
partial_product_22(370) <= '0';
partial_product_22(371) <= '0';
partial_product_22(372) <= '0';
partial_product_22(373) <= '0';
partial_product_22(374) <= '0';
partial_product_22(375) <= '0';
partial_product_22(376) <= '0';
partial_product_22(377) <= '0';
partial_product_22(378) <= '0';
partial_product_22(379) <= '0';
partial_product_22(380) <= '0';
partial_product_22(381) <= '0';
partial_product_22(382) <= '0';
partial_product_22(383) <= '0';
partial_product_22(384) <= '0';
partial_product_22(385) <= '0';
partial_product_22(386) <= '0';
partial_product_22(387) <= '0';
partial_product_22(388) <= '0';
partial_product_22(389) <= '0';
partial_product_22(390) <= '0';
partial_product_22(391) <= '0';
partial_product_22(392) <= '0';
partial_product_22(393) <= '0';
partial_product_22(394) <= '0';
partial_product_22(395) <= '0';
partial_product_22(396) <= '0';
partial_product_22(397) <= '0';
partial_product_22(398) <= '0';
partial_product_22(399) <= '0';
partial_product_22(400) <= '0';
partial_product_22(401) <= '0';
partial_product_22(402) <= '0';
partial_product_22(403) <= '0';
partial_product_22(404) <= '0';
partial_product_22(405) <= '0';
partial_product_22(406) <= '0';
partial_product_22(407) <= '0';
partial_product_22(408) <= '0';
partial_product_22(409) <= '0';
partial_product_22(410) <= '0';
partial_product_22(411) <= '0';
partial_product_22(412) <= '0';
partial_product_22(413) <= '0';
partial_product_22(414) <= '0';
partial_product_22(415) <= '0';
partial_product_22(416) <= '0';
partial_product_22(417) <= '0';
partial_product_22(418) <= '0';
partial_product_22(419) <= '0';
partial_product_22(420) <= '0';
partial_product_22(421) <= '0';
partial_product_22(422) <= '0';
partial_product_22(423) <= '0';
partial_product_22(424) <= '0';
partial_product_22(425) <= '0';
partial_product_22(426) <= '0';
partial_product_22(427) <= '0';
partial_product_22(428) <= '0';
partial_product_22(429) <= '0';
partial_product_22(430) <= '0';
partial_product_22(431) <= '0';
partial_product_22(432) <= '0';
partial_product_22(433) <= '0';
partial_product_22(434) <= '0';
partial_product_22(435) <= '0';
partial_product_22(436) <= '0';
partial_product_22(437) <= '0';
partial_product_22(438) <= '0';
partial_product_22(439) <= '0';
partial_product_22(440) <= '0';
partial_product_22(441) <= '0';
partial_product_22(442) <= '0';
partial_product_22(443) <= '0';
partial_product_22(444) <= '0';
partial_product_22(445) <= '0';
partial_product_22(446) <= '0';
partial_product_22(447) <= '0';
partial_product_22(448) <= '0';
partial_product_22(449) <= '0';
partial_product_22(450) <= '0';
partial_product_22(451) <= '0';
partial_product_22(452) <= '0';
partial_product_22(453) <= '0';
partial_product_22(454) <= '0';
partial_product_22(455) <= '0';
partial_product_22(456) <= '0';
partial_product_22(457) <= '0';
partial_product_22(458) <= '0';
partial_product_22(459) <= '0';
partial_product_22(460) <= '0';
partial_product_22(461) <= '0';
partial_product_22(462) <= '0';
partial_product_22(463) <= '0';
partial_product_22(464) <= '0';
partial_product_22(465) <= '0';
partial_product_22(466) <= '0';
partial_product_22(467) <= '0';
partial_product_22(468) <= '0';
partial_product_22(469) <= '0';
partial_product_22(470) <= '0';
partial_product_22(471) <= '0';
partial_product_22(472) <= '0';
partial_product_22(473) <= '0';
partial_product_22(474) <= '0';
partial_product_22(475) <= '0';
partial_product_22(476) <= '0';
partial_product_22(477) <= '0';
partial_product_22(478) <= '0';
partial_product_22(479) <= '0';
partial_product_22(480) <= '0';
partial_product_22(481) <= '0';
partial_product_22(482) <= '0';
partial_product_22(483) <= '0';
partial_product_22(484) <= '0';
partial_product_22(485) <= '0';
partial_product_22(486) <= '0';
partial_product_22(487) <= '0';
partial_product_22(488) <= '0';
partial_product_22(489) <= '0';
partial_product_22(490) <= '0';
partial_product_22(491) <= '0';
partial_product_22(492) <= '0';
partial_product_22(493) <= '0';
partial_product_22(494) <= '0';
partial_product_22(495) <= '0';
partial_product_22(496) <= '0';
partial_product_22(497) <= '0';
partial_product_22(498) <= '0';
partial_product_22(499) <= '0';
partial_product_22(500) <= '0';
partial_product_22(501) <= '0';
partial_product_22(502) <= '0';
partial_product_22(503) <= '0';
partial_product_22(504) <= '0';
partial_product_22(505) <= '0';
partial_product_22(506) <= '0';
partial_product_22(507) <= '0';
partial_product_22(508) <= '0';
partial_product_22(509) <= '0';
partial_product_22(510) <= '0';
partial_product_22(511) <= '0';
partial_product_22(512) <= '0';
partial_product_23(0) <= '0';
partial_product_23(1) <= '0';
partial_product_23(2) <= '0';
partial_product_23(3) <= '0';
partial_product_23(4) <= '0';
partial_product_23(5) <= '0';
partial_product_23(6) <= '0';
partial_product_23(7) <= '0';
partial_product_23(8) <= '0';
partial_product_23(9) <= '0';
partial_product_23(10) <= '0';
partial_product_23(11) <= '0';
partial_product_23(12) <= '0';
partial_product_23(13) <= '0';
partial_product_23(14) <= '0';
partial_product_23(15) <= '0';
partial_product_23(16) <= '0';
partial_product_23(17) <= '0';
partial_product_23(18) <= '0';
partial_product_23(19) <= '0';
partial_product_23(20) <= '0';
partial_product_23(21) <= '0';
partial_product_23(22) <= '0';
partial_product_23(23) <= '0';
partial_product_23(24) <= '0';
partial_product_23(25) <= '0';
partial_product_23(26) <= '0';
partial_product_23(27) <= '0';
partial_product_23(28) <= '0';
partial_product_23(29) <= '0';
partial_product_23(30) <= '0';
partial_product_23(31) <= '0';
partial_product_23(32) <= '0';
partial_product_23(33) <= '0';
partial_product_23(34) <= '0';
partial_product_23(35) <= '0';
partial_product_23(36) <= '0';
partial_product_23(37) <= '0';
partial_product_23(38) <= '0';
partial_product_23(39) <= '0';
partial_product_23(40) <= '0';
partial_product_23(41) <= '0';
partial_product_23(42) <= '0';
partial_product_23(43) <= '0';
partial_product_23(44) <= '0';
partial_product_23(45) <= '0';
partial_product_23(46) <= '0';
partial_product_23(47) <= '0';
partial_product_23(48) <= '0';
partial_product_23(49) <= '0';
partial_product_23(50) <= '0';
partial_product_23(51) <= '0';
partial_product_23(52) <= '0';
partial_product_23(53) <= '0';
partial_product_23(54) <= '0';
partial_product_23(55) <= '0';
partial_product_23(56) <= '0';
partial_product_23(57) <= '0';
partial_product_23(58) <= '0';
partial_product_23(59) <= '0';
partial_product_23(60) <= '0';
partial_product_23(61) <= '0';
partial_product_23(62) <= '0';
partial_product_23(63) <= '0';
partial_product_23(64) <= '0';
partial_product_23(65) <= '0';
partial_product_23(66) <= '0';
partial_product_23(67) <= '0';
partial_product_23(68) <= '0';
partial_product_23(69) <= '0';
partial_product_23(70) <= '0';
partial_product_23(71) <= '0';
partial_product_23(72) <= '0';
partial_product_23(73) <= '0';
partial_product_23(74) <= '0';
partial_product_23(75) <= '0';
partial_product_23(76) <= '0';
partial_product_23(77) <= '0';
partial_product_23(78) <= '0';
partial_product_23(79) <= '0';
partial_product_23(80) <= '0';
partial_product_23(81) <= '0';
partial_product_23(82) <= '0';
partial_product_23(83) <= '0';
partial_product_23(84) <= '0';
partial_product_23(85) <= '0';
partial_product_23(86) <= '0';
partial_product_23(87) <= '0';
partial_product_23(88) <= '0';
partial_product_23(89) <= '0';
partial_product_23(90) <= '0';
partial_product_23(91) <= '0';
partial_product_23(92) <= '0';
partial_product_23(93) <= '0';
partial_product_23(94) <= '0';
partial_product_23(95) <= '0';
partial_product_23(96) <= '0';
partial_product_23(97) <= '0';
partial_product_23(98) <= '0';
partial_product_23(99) <= '0';
partial_product_23(100) <= '0';
partial_product_23(101) <= '0';
partial_product_23(102) <= '0';
partial_product_23(103) <= '0';
partial_product_23(104) <= '0';
partial_product_23(105) <= '0';
partial_product_23(106) <= '0';
partial_product_23(107) <= '0';
partial_product_23(108) <= '0';
partial_product_23(109) <= '0';
partial_product_23(110) <= '0';
partial_product_23(111) <= '0';
partial_product_23(112) <= '0';
partial_product_23(113) <= '0';
partial_product_23(114) <= '0';
partial_product_23(115) <= '0';
partial_product_23(116) <= '0';
partial_product_23(117) <= '0';
partial_product_23(118) <= '0';
partial_product_23(119) <= '0';
partial_product_23(120) <= '0';
partial_product_23(121) <= '0';
partial_product_23(122) <= '0';
partial_product_23(123) <= '0';
partial_product_23(124) <= '0';
partial_product_23(125) <= '0';
partial_product_23(126) <= '0';
partial_product_23(127) <= '0';
partial_product_23(128) <= '0';
partial_product_23(129) <= '0';
partial_product_23(130) <= '0';
partial_product_23(131) <= '0';
partial_product_23(132) <= '0';
partial_product_23(133) <= '0';
partial_product_23(134) <= '0';
partial_product_23(135) <= '0';
partial_product_23(136) <= '0';
partial_product_23(137) <= '0';
partial_product_23(138) <= '0';
partial_product_23(139) <= '0';
partial_product_23(140) <= '0';
partial_product_23(141) <= '0';
partial_product_23(142) <= '0';
partial_product_23(143) <= '0';
partial_product_23(144) <= '0';
partial_product_23(145) <= '0';
partial_product_23(146) <= '0';
partial_product_23(147) <= '0';
partial_product_23(148) <= '0';
partial_product_23(149) <= '0';
partial_product_23(150) <= '0';
partial_product_23(151) <= '0';
partial_product_23(152) <= '0';
partial_product_23(153) <= '0';
partial_product_23(154) <= '0';
partial_product_23(155) <= '0';
partial_product_23(156) <= '0';
partial_product_23(157) <= '0';
partial_product_23(158) <= '0';
partial_product_23(159) <= '0';
partial_product_23(160) <= '0';
partial_product_23(161) <= '0';
partial_product_23(162) <= '0';
partial_product_23(163) <= '0';
partial_product_23(164) <= '0';
partial_product_23(165) <= '0';
partial_product_23(166) <= '0';
partial_product_23(167) <= '0';
partial_product_23(168) <= '0';
partial_product_23(169) <= '0';
partial_product_23(170) <= '0';
partial_product_23(171) <= '0';
partial_product_23(172) <= '0';
partial_product_23(173) <= '0';
partial_product_23(174) <= '0';
partial_product_23(175) <= '0';
partial_product_23(176) <= '0';
partial_product_23(177) <= '0';
partial_product_23(178) <= '0';
partial_product_23(179) <= '0';
partial_product_23(180) <= '0';
partial_product_23(181) <= '0';
partial_product_23(182) <= '0';
partial_product_23(183) <= '0';
partial_product_23(184) <= '0';
partial_product_23(185) <= '0';
partial_product_23(186) <= '0';
partial_product_23(187) <= '0';
partial_product_23(188) <= '0';
partial_product_23(189) <= '0';
partial_product_23(190) <= '0';
partial_product_23(191) <= '0';
partial_product_23(192) <= '0';
partial_product_23(193) <= '0';
partial_product_23(194) <= '0';
partial_product_23(195) <= '0';
partial_product_23(196) <= '0';
partial_product_23(197) <= '0';
partial_product_23(198) <= '0';
partial_product_23(199) <= '0';
partial_product_23(200) <= '0';
partial_product_23(201) <= '0';
partial_product_23(202) <= '0';
partial_product_23(203) <= '0';
partial_product_23(204) <= '0';
partial_product_23(205) <= '0';
partial_product_23(206) <= '0';
partial_product_23(207) <= '0';
partial_product_23(208) <= '0';
partial_product_23(209) <= '0';
partial_product_23(210) <= '0';
partial_product_23(211) <= '0';
partial_product_23(212) <= '0';
partial_product_23(213) <= '0';
partial_product_23(214) <= '0';
partial_product_23(215) <= '0';
partial_product_23(216) <= '0';
partial_product_23(217) <= '0';
partial_product_23(218) <= '0';
partial_product_23(219) <= '0';
partial_product_23(220) <= '0';
partial_product_23(221) <= '0';
partial_product_23(222) <= '0';
partial_product_23(223) <= '0';
partial_product_23(224) <= '0';
partial_product_23(225) <= '0';
partial_product_23(226) <= '0';
partial_product_23(227) <= '0';
partial_product_23(228) <= '0';
partial_product_23(229) <= '0';
partial_product_23(230) <= '0';
partial_product_23(231) <= '0';
partial_product_23(232) <= '0';
partial_product_23(233) <= '0';
partial_product_23(234) <= '0';
partial_product_23(235) <= '0';
partial_product_23(236) <= '0';
partial_product_23(237) <= '0';
partial_product_23(238) <= temp_mult_86(238);
partial_product_23(239) <= temp_mult_86(239);
partial_product_23(240) <= temp_mult_86(240);
partial_product_23(241) <= temp_mult_86(241);
partial_product_23(242) <= temp_mult_86(242);
partial_product_23(243) <= temp_mult_86(243);
partial_product_23(244) <= temp_mult_86(244);
partial_product_23(245) <= temp_mult_86(245);
partial_product_23(246) <= temp_mult_86(246);
partial_product_23(247) <= temp_mult_86(247);
partial_product_23(248) <= temp_mult_86(248);
partial_product_23(249) <= temp_mult_86(249);
partial_product_23(250) <= temp_mult_86(250);
partial_product_23(251) <= temp_mult_86(251);
partial_product_23(252) <= temp_mult_86(252);
partial_product_23(253) <= temp_mult_86(253);
partial_product_23(254) <= temp_mult_86(254);
partial_product_23(255) <= temp_mult_86(255);
partial_product_23(256) <= temp_mult_86(256);
partial_product_23(257) <= temp_mult_86(257);
partial_product_23(258) <= temp_mult_86(258);
partial_product_23(259) <= temp_mult_86(259);
partial_product_23(260) <= temp_mult_86(260);
partial_product_23(261) <= temp_mult_86(261);
partial_product_23(262) <= temp_mult_86(262);
partial_product_23(263) <= temp_mult_86(263);
partial_product_23(264) <= temp_mult_86(264);
partial_product_23(265) <= temp_mult_86(265);
partial_product_23(266) <= temp_mult_86(266);
partial_product_23(267) <= temp_mult_86(267);
partial_product_23(268) <= temp_mult_86(268);
partial_product_23(269) <= temp_mult_86(269);
partial_product_23(270) <= temp_mult_86(270);
partial_product_23(271) <= temp_mult_86(271);
partial_product_23(272) <= temp_mult_86(272);
partial_product_23(273) <= temp_mult_86(273);
partial_product_23(274) <= temp_mult_86(274);
partial_product_23(275) <= temp_mult_86(275);
partial_product_23(276) <= temp_mult_86(276);
partial_product_23(277) <= temp_mult_86(277);
partial_product_23(278) <= temp_mult_86(278);
partial_product_23(279) <= '0';
partial_product_23(280) <= '0';
partial_product_23(281) <= '0';
partial_product_23(282) <= '0';
partial_product_23(283) <= '0';
partial_product_23(284) <= '0';
partial_product_23(285) <= '0';
partial_product_23(286) <= '0';
partial_product_23(287) <= '0';
partial_product_23(288) <= '0';
partial_product_23(289) <= '0';
partial_product_23(290) <= '0';
partial_product_23(291) <= '0';
partial_product_23(292) <= '0';
partial_product_23(293) <= '0';
partial_product_23(294) <= '0';
partial_product_23(295) <= '0';
partial_product_23(296) <= '0';
partial_product_23(297) <= '0';
partial_product_23(298) <= '0';
partial_product_23(299) <= '0';
partial_product_23(300) <= '0';
partial_product_23(301) <= '0';
partial_product_23(302) <= '0';
partial_product_23(303) <= '0';
partial_product_23(304) <= '0';
partial_product_23(305) <= '0';
partial_product_23(306) <= '0';
partial_product_23(307) <= '0';
partial_product_23(308) <= '0';
partial_product_23(309) <= '0';
partial_product_23(310) <= '0';
partial_product_23(311) <= '0';
partial_product_23(312) <= '0';
partial_product_23(313) <= '0';
partial_product_23(314) <= '0';
partial_product_23(315) <= '0';
partial_product_23(316) <= '0';
partial_product_23(317) <= '0';
partial_product_23(318) <= '0';
partial_product_23(319) <= '0';
partial_product_23(320) <= '0';
partial_product_23(321) <= '0';
partial_product_23(322) <= '0';
partial_product_23(323) <= '0';
partial_product_23(324) <= '0';
partial_product_23(325) <= '0';
partial_product_23(326) <= '0';
partial_product_23(327) <= '0';
partial_product_23(328) <= '0';
partial_product_23(329) <= '0';
partial_product_23(330) <= '0';
partial_product_23(331) <= '0';
partial_product_23(332) <= '0';
partial_product_23(333) <= '0';
partial_product_23(334) <= '0';
partial_product_23(335) <= '0';
partial_product_23(336) <= '0';
partial_product_23(337) <= '0';
partial_product_23(338) <= '0';
partial_product_23(339) <= '0';
partial_product_23(340) <= '0';
partial_product_23(341) <= '0';
partial_product_23(342) <= '0';
partial_product_23(343) <= '0';
partial_product_23(344) <= '0';
partial_product_23(345) <= '0';
partial_product_23(346) <= '0';
partial_product_23(347) <= '0';
partial_product_23(348) <= '0';
partial_product_23(349) <= '0';
partial_product_23(350) <= '0';
partial_product_23(351) <= '0';
partial_product_23(352) <= '0';
partial_product_23(353) <= '0';
partial_product_23(354) <= '0';
partial_product_23(355) <= '0';
partial_product_23(356) <= '0';
partial_product_23(357) <= '0';
partial_product_23(358) <= '0';
partial_product_23(359) <= '0';
partial_product_23(360) <= '0';
partial_product_23(361) <= '0';
partial_product_23(362) <= '0';
partial_product_23(363) <= '0';
partial_product_23(364) <= '0';
partial_product_23(365) <= '0';
partial_product_23(366) <= '0';
partial_product_23(367) <= '0';
partial_product_23(368) <= '0';
partial_product_23(369) <= '0';
partial_product_23(370) <= '0';
partial_product_23(371) <= '0';
partial_product_23(372) <= '0';
partial_product_23(373) <= '0';
partial_product_23(374) <= '0';
partial_product_23(375) <= '0';
partial_product_23(376) <= '0';
partial_product_23(377) <= '0';
partial_product_23(378) <= '0';
partial_product_23(379) <= '0';
partial_product_23(380) <= '0';
partial_product_23(381) <= '0';
partial_product_23(382) <= '0';
partial_product_23(383) <= '0';
partial_product_23(384) <= '0';
partial_product_23(385) <= '0';
partial_product_23(386) <= '0';
partial_product_23(387) <= '0';
partial_product_23(388) <= '0';
partial_product_23(389) <= '0';
partial_product_23(390) <= '0';
partial_product_23(391) <= '0';
partial_product_23(392) <= '0';
partial_product_23(393) <= '0';
partial_product_23(394) <= '0';
partial_product_23(395) <= '0';
partial_product_23(396) <= '0';
partial_product_23(397) <= '0';
partial_product_23(398) <= '0';
partial_product_23(399) <= '0';
partial_product_23(400) <= '0';
partial_product_23(401) <= '0';
partial_product_23(402) <= '0';
partial_product_23(403) <= '0';
partial_product_23(404) <= '0';
partial_product_23(405) <= '0';
partial_product_23(406) <= '0';
partial_product_23(407) <= '0';
partial_product_23(408) <= '0';
partial_product_23(409) <= '0';
partial_product_23(410) <= '0';
partial_product_23(411) <= '0';
partial_product_23(412) <= '0';
partial_product_23(413) <= '0';
partial_product_23(414) <= '0';
partial_product_23(415) <= '0';
partial_product_23(416) <= '0';
partial_product_23(417) <= '0';
partial_product_23(418) <= '0';
partial_product_23(419) <= '0';
partial_product_23(420) <= '0';
partial_product_23(421) <= '0';
partial_product_23(422) <= '0';
partial_product_23(423) <= '0';
partial_product_23(424) <= '0';
partial_product_23(425) <= '0';
partial_product_23(426) <= '0';
partial_product_23(427) <= '0';
partial_product_23(428) <= '0';
partial_product_23(429) <= '0';
partial_product_23(430) <= '0';
partial_product_23(431) <= '0';
partial_product_23(432) <= '0';
partial_product_23(433) <= '0';
partial_product_23(434) <= '0';
partial_product_23(435) <= '0';
partial_product_23(436) <= '0';
partial_product_23(437) <= '0';
partial_product_23(438) <= '0';
partial_product_23(439) <= '0';
partial_product_23(440) <= '0';
partial_product_23(441) <= '0';
partial_product_23(442) <= '0';
partial_product_23(443) <= '0';
partial_product_23(444) <= '0';
partial_product_23(445) <= '0';
partial_product_23(446) <= '0';
partial_product_23(447) <= '0';
partial_product_23(448) <= '0';
partial_product_23(449) <= '0';
partial_product_23(450) <= '0';
partial_product_23(451) <= '0';
partial_product_23(452) <= '0';
partial_product_23(453) <= '0';
partial_product_23(454) <= '0';
partial_product_23(455) <= '0';
partial_product_23(456) <= '0';
partial_product_23(457) <= '0';
partial_product_23(458) <= '0';
partial_product_23(459) <= '0';
partial_product_23(460) <= '0';
partial_product_23(461) <= '0';
partial_product_23(462) <= '0';
partial_product_23(463) <= '0';
partial_product_23(464) <= '0';
partial_product_23(465) <= '0';
partial_product_23(466) <= '0';
partial_product_23(467) <= '0';
partial_product_23(468) <= '0';
partial_product_23(469) <= '0';
partial_product_23(470) <= '0';
partial_product_23(471) <= '0';
partial_product_23(472) <= '0';
partial_product_23(473) <= '0';
partial_product_23(474) <= '0';
partial_product_23(475) <= '0';
partial_product_23(476) <= '0';
partial_product_23(477) <= '0';
partial_product_23(478) <= '0';
partial_product_23(479) <= '0';
partial_product_23(480) <= '0';
partial_product_23(481) <= '0';
partial_product_23(482) <= '0';
partial_product_23(483) <= '0';
partial_product_23(484) <= '0';
partial_product_23(485) <= '0';
partial_product_23(486) <= '0';
partial_product_23(487) <= '0';
partial_product_23(488) <= '0';
partial_product_23(489) <= '0';
partial_product_23(490) <= '0';
partial_product_23(491) <= '0';
partial_product_23(492) <= '0';
partial_product_23(493) <= '0';
partial_product_23(494) <= '0';
partial_product_23(495) <= '0';
partial_product_23(496) <= '0';
partial_product_23(497) <= '0';
partial_product_23(498) <= '0';
partial_product_23(499) <= '0';
partial_product_23(500) <= '0';
partial_product_23(501) <= '0';
partial_product_23(502) <= '0';
partial_product_23(503) <= '0';
partial_product_23(504) <= '0';
partial_product_23(505) <= '0';
partial_product_23(506) <= '0';
partial_product_23(507) <= '0';
partial_product_23(508) <= '0';
partial_product_23(509) <= '0';
partial_product_23(510) <= '0';
partial_product_23(511) <= '0';
partial_product_23(512) <= '0';
partial_product_24(0) <= '0';
partial_product_24(1) <= '0';
partial_product_24(2) <= '0';
partial_product_24(3) <= '0';
partial_product_24(4) <= '0';
partial_product_24(5) <= '0';
partial_product_24(6) <= '0';
partial_product_24(7) <= '0';
partial_product_24(8) <= '0';
partial_product_24(9) <= '0';
partial_product_24(10) <= '0';
partial_product_24(11) <= '0';
partial_product_24(12) <= '0';
partial_product_24(13) <= '0';
partial_product_24(14) <= '0';
partial_product_24(15) <= '0';
partial_product_24(16) <= '0';
partial_product_24(17) <= '0';
partial_product_24(18) <= '0';
partial_product_24(19) <= '0';
partial_product_24(20) <= '0';
partial_product_24(21) <= '0';
partial_product_24(22) <= '0';
partial_product_24(23) <= '0';
partial_product_24(24) <= '0';
partial_product_24(25) <= '0';
partial_product_24(26) <= '0';
partial_product_24(27) <= '0';
partial_product_24(28) <= '0';
partial_product_24(29) <= '0';
partial_product_24(30) <= '0';
partial_product_24(31) <= '0';
partial_product_24(32) <= '0';
partial_product_24(33) <= '0';
partial_product_24(34) <= '0';
partial_product_24(35) <= '0';
partial_product_24(36) <= '0';
partial_product_24(37) <= '0';
partial_product_24(38) <= '0';
partial_product_24(39) <= '0';
partial_product_24(40) <= '0';
partial_product_24(41) <= '0';
partial_product_24(42) <= '0';
partial_product_24(43) <= '0';
partial_product_24(44) <= '0';
partial_product_24(45) <= '0';
partial_product_24(46) <= '0';
partial_product_24(47) <= '0';
partial_product_24(48) <= '0';
partial_product_24(49) <= '0';
partial_product_24(50) <= '0';
partial_product_24(51) <= '0';
partial_product_24(52) <= '0';
partial_product_24(53) <= '0';
partial_product_24(54) <= '0';
partial_product_24(55) <= '0';
partial_product_24(56) <= '0';
partial_product_24(57) <= '0';
partial_product_24(58) <= '0';
partial_product_24(59) <= '0';
partial_product_24(60) <= '0';
partial_product_24(61) <= '0';
partial_product_24(62) <= '0';
partial_product_24(63) <= '0';
partial_product_24(64) <= '0';
partial_product_24(65) <= '0';
partial_product_24(66) <= '0';
partial_product_24(67) <= '0';
partial_product_24(68) <= '0';
partial_product_24(69) <= '0';
partial_product_24(70) <= '0';
partial_product_24(71) <= '0';
partial_product_24(72) <= '0';
partial_product_24(73) <= '0';
partial_product_24(74) <= '0';
partial_product_24(75) <= '0';
partial_product_24(76) <= '0';
partial_product_24(77) <= '0';
partial_product_24(78) <= '0';
partial_product_24(79) <= '0';
partial_product_24(80) <= '0';
partial_product_24(81) <= '0';
partial_product_24(82) <= '0';
partial_product_24(83) <= '0';
partial_product_24(84) <= '0';
partial_product_24(85) <= '0';
partial_product_24(86) <= '0';
partial_product_24(87) <= '0';
partial_product_24(88) <= '0';
partial_product_24(89) <= '0';
partial_product_24(90) <= '0';
partial_product_24(91) <= '0';
partial_product_24(92) <= '0';
partial_product_24(93) <= '0';
partial_product_24(94) <= '0';
partial_product_24(95) <= '0';
partial_product_24(96) <= '0';
partial_product_24(97) <= '0';
partial_product_24(98) <= '0';
partial_product_24(99) <= '0';
partial_product_24(100) <= '0';
partial_product_24(101) <= '0';
partial_product_24(102) <= '0';
partial_product_24(103) <= '0';
partial_product_24(104) <= '0';
partial_product_24(105) <= '0';
partial_product_24(106) <= '0';
partial_product_24(107) <= '0';
partial_product_24(108) <= '0';
partial_product_24(109) <= '0';
partial_product_24(110) <= '0';
partial_product_24(111) <= '0';
partial_product_24(112) <= '0';
partial_product_24(113) <= '0';
partial_product_24(114) <= '0';
partial_product_24(115) <= '0';
partial_product_24(116) <= '0';
partial_product_24(117) <= '0';
partial_product_24(118) <= '0';
partial_product_24(119) <= '0';
partial_product_24(120) <= '0';
partial_product_24(121) <= '0';
partial_product_24(122) <= '0';
partial_product_24(123) <= '0';
partial_product_24(124) <= '0';
partial_product_24(125) <= '0';
partial_product_24(126) <= '0';
partial_product_24(127) <= '0';
partial_product_24(128) <= '0';
partial_product_24(129) <= '0';
partial_product_24(130) <= '0';
partial_product_24(131) <= '0';
partial_product_24(132) <= '0';
partial_product_24(133) <= '0';
partial_product_24(134) <= '0';
partial_product_24(135) <= '0';
partial_product_24(136) <= '0';
partial_product_24(137) <= '0';
partial_product_24(138) <= '0';
partial_product_24(139) <= '0';
partial_product_24(140) <= '0';
partial_product_24(141) <= '0';
partial_product_24(142) <= '0';
partial_product_24(143) <= '0';
partial_product_24(144) <= '0';
partial_product_24(145) <= '0';
partial_product_24(146) <= '0';
partial_product_24(147) <= '0';
partial_product_24(148) <= '0';
partial_product_24(149) <= '0';
partial_product_24(150) <= '0';
partial_product_24(151) <= '0';
partial_product_24(152) <= '0';
partial_product_24(153) <= '0';
partial_product_24(154) <= '0';
partial_product_24(155) <= '0';
partial_product_24(156) <= '0';
partial_product_24(157) <= '0';
partial_product_24(158) <= '0';
partial_product_24(159) <= '0';
partial_product_24(160) <= '0';
partial_product_24(161) <= '0';
partial_product_24(162) <= '0';
partial_product_24(163) <= '0';
partial_product_24(164) <= '0';
partial_product_24(165) <= '0';
partial_product_24(166) <= '0';
partial_product_24(167) <= '0';
partial_product_24(168) <= '0';
partial_product_24(169) <= '0';
partial_product_24(170) <= '0';
partial_product_24(171) <= '0';
partial_product_24(172) <= '0';
partial_product_24(173) <= '0';
partial_product_24(174) <= '0';
partial_product_24(175) <= '0';
partial_product_24(176) <= '0';
partial_product_24(177) <= '0';
partial_product_24(178) <= '0';
partial_product_24(179) <= '0';
partial_product_24(180) <= '0';
partial_product_24(181) <= '0';
partial_product_24(182) <= '0';
partial_product_24(183) <= '0';
partial_product_24(184) <= '0';
partial_product_24(185) <= '0';
partial_product_24(186) <= '0';
partial_product_24(187) <= '0';
partial_product_24(188) <= '0';
partial_product_24(189) <= '0';
partial_product_24(190) <= '0';
partial_product_24(191) <= '0';
partial_product_24(192) <= '0';
partial_product_24(193) <= '0';
partial_product_24(194) <= '0';
partial_product_24(195) <= '0';
partial_product_24(196) <= '0';
partial_product_24(197) <= '0';
partial_product_24(198) <= '0';
partial_product_24(199) <= '0';
partial_product_24(200) <= '0';
partial_product_24(201) <= '0';
partial_product_24(202) <= '0';
partial_product_24(203) <= '0';
partial_product_24(204) <= '0';
partial_product_24(205) <= '0';
partial_product_24(206) <= '0';
partial_product_24(207) <= '0';
partial_product_24(208) <= '0';
partial_product_24(209) <= '0';
partial_product_24(210) <= '0';
partial_product_24(211) <= '0';
partial_product_24(212) <= '0';
partial_product_24(213) <= '0';
partial_product_24(214) <= '0';
partial_product_24(215) <= '0';
partial_product_24(216) <= '0';
partial_product_24(217) <= '0';
partial_product_24(218) <= '0';
partial_product_24(219) <= '0';
partial_product_24(220) <= '0';
partial_product_24(221) <= '0';
partial_product_24(222) <= '0';
partial_product_24(223) <= '0';
partial_product_24(224) <= '0';
partial_product_24(225) <= '0';
partial_product_24(226) <= '0';
partial_product_24(227) <= '0';
partial_product_24(228) <= '0';
partial_product_24(229) <= '0';
partial_product_24(230) <= '0';
partial_product_24(231) <= '0';
partial_product_24(232) <= '0';
partial_product_24(233) <= '0';
partial_product_24(234) <= '0';
partial_product_24(235) <= '0';
partial_product_24(236) <= '0';
partial_product_24(237) <= '0';
partial_product_24(238) <= '0';
partial_product_24(239) <= '0';
partial_product_24(240) <= temp_mult_160(240);
partial_product_24(241) <= temp_mult_160(241);
partial_product_24(242) <= temp_mult_160(242);
partial_product_24(243) <= temp_mult_160(243);
partial_product_24(244) <= temp_mult_160(244);
partial_product_24(245) <= temp_mult_160(245);
partial_product_24(246) <= temp_mult_160(246);
partial_product_24(247) <= temp_mult_160(247);
partial_product_24(248) <= temp_mult_160(248);
partial_product_24(249) <= temp_mult_160(249);
partial_product_24(250) <= temp_mult_160(250);
partial_product_24(251) <= temp_mult_160(251);
partial_product_24(252) <= temp_mult_160(252);
partial_product_24(253) <= temp_mult_160(253);
partial_product_24(254) <= temp_mult_160(254);
partial_product_24(255) <= temp_mult_160(255);
partial_product_24(256) <= temp_mult_160(256);
partial_product_24(257) <= temp_mult_160(257);
partial_product_24(258) <= temp_mult_160(258);
partial_product_24(259) <= temp_mult_160(259);
partial_product_24(260) <= temp_mult_160(260);
partial_product_24(261) <= temp_mult_160(261);
partial_product_24(262) <= temp_mult_160(262);
partial_product_24(263) <= temp_mult_160(263);
partial_product_24(264) <= temp_mult_160(264);
partial_product_24(265) <= temp_mult_160(265);
partial_product_24(266) <= temp_mult_160(266);
partial_product_24(267) <= temp_mult_160(267);
partial_product_24(268) <= temp_mult_160(268);
partial_product_24(269) <= temp_mult_160(269);
partial_product_24(270) <= temp_mult_160(270);
partial_product_24(271) <= temp_mult_160(271);
partial_product_24(272) <= '0';
partial_product_24(273) <= '0';
partial_product_24(274) <= '0';
partial_product_24(275) <= '0';
partial_product_24(276) <= '0';
partial_product_24(277) <= '0';
partial_product_24(278) <= '0';
partial_product_24(279) <= '0';
partial_product_24(280) <= '0';
partial_product_24(281) <= '0';
partial_product_24(282) <= '0';
partial_product_24(283) <= '0';
partial_product_24(284) <= '0';
partial_product_24(285) <= '0';
partial_product_24(286) <= '0';
partial_product_24(287) <= '0';
partial_product_24(288) <= '0';
partial_product_24(289) <= '0';
partial_product_24(290) <= '0';
partial_product_24(291) <= '0';
partial_product_24(292) <= '0';
partial_product_24(293) <= '0';
partial_product_24(294) <= '0';
partial_product_24(295) <= '0';
partial_product_24(296) <= '0';
partial_product_24(297) <= '0';
partial_product_24(298) <= '0';
partial_product_24(299) <= '0';
partial_product_24(300) <= '0';
partial_product_24(301) <= '0';
partial_product_24(302) <= '0';
partial_product_24(303) <= '0';
partial_product_24(304) <= '0';
partial_product_24(305) <= '0';
partial_product_24(306) <= '0';
partial_product_24(307) <= '0';
partial_product_24(308) <= '0';
partial_product_24(309) <= '0';
partial_product_24(310) <= '0';
partial_product_24(311) <= '0';
partial_product_24(312) <= '0';
partial_product_24(313) <= '0';
partial_product_24(314) <= '0';
partial_product_24(315) <= '0';
partial_product_24(316) <= '0';
partial_product_24(317) <= '0';
partial_product_24(318) <= '0';
partial_product_24(319) <= '0';
partial_product_24(320) <= '0';
partial_product_24(321) <= '0';
partial_product_24(322) <= '0';
partial_product_24(323) <= '0';
partial_product_24(324) <= '0';
partial_product_24(325) <= '0';
partial_product_24(326) <= '0';
partial_product_24(327) <= '0';
partial_product_24(328) <= '0';
partial_product_24(329) <= '0';
partial_product_24(330) <= '0';
partial_product_24(331) <= '0';
partial_product_24(332) <= '0';
partial_product_24(333) <= '0';
partial_product_24(334) <= '0';
partial_product_24(335) <= '0';
partial_product_24(336) <= '0';
partial_product_24(337) <= '0';
partial_product_24(338) <= '0';
partial_product_24(339) <= '0';
partial_product_24(340) <= '0';
partial_product_24(341) <= '0';
partial_product_24(342) <= '0';
partial_product_24(343) <= '0';
partial_product_24(344) <= '0';
partial_product_24(345) <= '0';
partial_product_24(346) <= '0';
partial_product_24(347) <= '0';
partial_product_24(348) <= '0';
partial_product_24(349) <= '0';
partial_product_24(350) <= '0';
partial_product_24(351) <= '0';
partial_product_24(352) <= '0';
partial_product_24(353) <= '0';
partial_product_24(354) <= '0';
partial_product_24(355) <= '0';
partial_product_24(356) <= '0';
partial_product_24(357) <= '0';
partial_product_24(358) <= '0';
partial_product_24(359) <= '0';
partial_product_24(360) <= '0';
partial_product_24(361) <= '0';
partial_product_24(362) <= '0';
partial_product_24(363) <= '0';
partial_product_24(364) <= '0';
partial_product_24(365) <= '0';
partial_product_24(366) <= '0';
partial_product_24(367) <= '0';
partial_product_24(368) <= '0';
partial_product_24(369) <= '0';
partial_product_24(370) <= '0';
partial_product_24(371) <= '0';
partial_product_24(372) <= '0';
partial_product_24(373) <= '0';
partial_product_24(374) <= '0';
partial_product_24(375) <= '0';
partial_product_24(376) <= '0';
partial_product_24(377) <= '0';
partial_product_24(378) <= '0';
partial_product_24(379) <= '0';
partial_product_24(380) <= '0';
partial_product_24(381) <= '0';
partial_product_24(382) <= '0';
partial_product_24(383) <= '0';
partial_product_24(384) <= '0';
partial_product_24(385) <= '0';
partial_product_24(386) <= '0';
partial_product_24(387) <= '0';
partial_product_24(388) <= '0';
partial_product_24(389) <= '0';
partial_product_24(390) <= '0';
partial_product_24(391) <= '0';
partial_product_24(392) <= '0';
partial_product_24(393) <= '0';
partial_product_24(394) <= '0';
partial_product_24(395) <= '0';
partial_product_24(396) <= '0';
partial_product_24(397) <= '0';
partial_product_24(398) <= '0';
partial_product_24(399) <= '0';
partial_product_24(400) <= '0';
partial_product_24(401) <= '0';
partial_product_24(402) <= '0';
partial_product_24(403) <= '0';
partial_product_24(404) <= '0';
partial_product_24(405) <= '0';
partial_product_24(406) <= '0';
partial_product_24(407) <= '0';
partial_product_24(408) <= '0';
partial_product_24(409) <= '0';
partial_product_24(410) <= '0';
partial_product_24(411) <= '0';
partial_product_24(412) <= '0';
partial_product_24(413) <= '0';
partial_product_24(414) <= '0';
partial_product_24(415) <= '0';
partial_product_24(416) <= '0';
partial_product_24(417) <= '0';
partial_product_24(418) <= '0';
partial_product_24(419) <= '0';
partial_product_24(420) <= '0';
partial_product_24(421) <= '0';
partial_product_24(422) <= '0';
partial_product_24(423) <= '0';
partial_product_24(424) <= '0';
partial_product_24(425) <= '0';
partial_product_24(426) <= '0';
partial_product_24(427) <= '0';
partial_product_24(428) <= '0';
partial_product_24(429) <= '0';
partial_product_24(430) <= '0';
partial_product_24(431) <= '0';
partial_product_24(432) <= '0';
partial_product_24(433) <= '0';
partial_product_24(434) <= '0';
partial_product_24(435) <= '0';
partial_product_24(436) <= '0';
partial_product_24(437) <= '0';
partial_product_24(438) <= '0';
partial_product_24(439) <= '0';
partial_product_24(440) <= '0';
partial_product_24(441) <= '0';
partial_product_24(442) <= '0';
partial_product_24(443) <= '0';
partial_product_24(444) <= '0';
partial_product_24(445) <= '0';
partial_product_24(446) <= '0';
partial_product_24(447) <= '0';
partial_product_24(448) <= '0';
partial_product_24(449) <= '0';
partial_product_24(450) <= '0';
partial_product_24(451) <= '0';
partial_product_24(452) <= '0';
partial_product_24(453) <= '0';
partial_product_24(454) <= '0';
partial_product_24(455) <= '0';
partial_product_24(456) <= '0';
partial_product_24(457) <= '0';
partial_product_24(458) <= '0';
partial_product_24(459) <= '0';
partial_product_24(460) <= '0';
partial_product_24(461) <= '0';
partial_product_24(462) <= '0';
partial_product_24(463) <= '0';
partial_product_24(464) <= '0';
partial_product_24(465) <= '0';
partial_product_24(466) <= '0';
partial_product_24(467) <= '0';
partial_product_24(468) <= '0';
partial_product_24(469) <= '0';
partial_product_24(470) <= '0';
partial_product_24(471) <= '0';
partial_product_24(472) <= '0';
partial_product_24(473) <= '0';
partial_product_24(474) <= '0';
partial_product_24(475) <= '0';
partial_product_24(476) <= '0';
partial_product_24(477) <= '0';
partial_product_24(478) <= '0';
partial_product_24(479) <= '0';
partial_product_24(480) <= '0';
partial_product_24(481) <= '0';
partial_product_24(482) <= '0';
partial_product_24(483) <= '0';
partial_product_24(484) <= '0';
partial_product_24(485) <= '0';
partial_product_24(486) <= '0';
partial_product_24(487) <= '0';
partial_product_24(488) <= '0';
partial_product_24(489) <= '0';
partial_product_24(490) <= '0';
partial_product_24(491) <= '0';
partial_product_24(492) <= '0';
partial_product_24(493) <= '0';
partial_product_24(494) <= '0';
partial_product_24(495) <= '0';
partial_product_24(496) <= '0';
partial_product_24(497) <= '0';
partial_product_24(498) <= '0';
partial_product_24(499) <= '0';
partial_product_24(500) <= '0';
partial_product_24(501) <= '0';
partial_product_24(502) <= '0';
partial_product_24(503) <= '0';
partial_product_24(504) <= '0';
partial_product_24(505) <= '0';
partial_product_24(506) <= '0';
partial_product_24(507) <= '0';
partial_product_24(508) <= '0';
partial_product_24(509) <= '0';
partial_product_24(510) <= '0';
partial_product_24(511) <= '0';
partial_product_24(512) <= '0';
partial_product_25(0) <= '0';
partial_product_25(1) <= '0';
partial_product_25(2) <= '0';
partial_product_25(3) <= '0';
partial_product_25(4) <= '0';
partial_product_25(5) <= '0';
partial_product_25(6) <= '0';
partial_product_25(7) <= '0';
partial_product_25(8) <= '0';
partial_product_25(9) <= '0';
partial_product_25(10) <= '0';
partial_product_25(11) <= '0';
partial_product_25(12) <= '0';
partial_product_25(13) <= '0';
partial_product_25(14) <= '0';
partial_product_25(15) <= '0';
partial_product_25(16) <= '0';
partial_product_25(17) <= '0';
partial_product_25(18) <= '0';
partial_product_25(19) <= '0';
partial_product_25(20) <= '0';
partial_product_25(21) <= '0';
partial_product_25(22) <= '0';
partial_product_25(23) <= '0';
partial_product_25(24) <= '0';
partial_product_25(25) <= '0';
partial_product_25(26) <= '0';
partial_product_25(27) <= '0';
partial_product_25(28) <= '0';
partial_product_25(29) <= '0';
partial_product_25(30) <= '0';
partial_product_25(31) <= '0';
partial_product_25(32) <= '0';
partial_product_25(33) <= '0';
partial_product_25(34) <= '0';
partial_product_25(35) <= '0';
partial_product_25(36) <= '0';
partial_product_25(37) <= '0';
partial_product_25(38) <= '0';
partial_product_25(39) <= '0';
partial_product_25(40) <= '0';
partial_product_25(41) <= '0';
partial_product_25(42) <= '0';
partial_product_25(43) <= '0';
partial_product_25(44) <= '0';
partial_product_25(45) <= '0';
partial_product_25(46) <= '0';
partial_product_25(47) <= '0';
partial_product_25(48) <= '0';
partial_product_25(49) <= '0';
partial_product_25(50) <= '0';
partial_product_25(51) <= '0';
partial_product_25(52) <= '0';
partial_product_25(53) <= '0';
partial_product_25(54) <= '0';
partial_product_25(55) <= '0';
partial_product_25(56) <= '0';
partial_product_25(57) <= '0';
partial_product_25(58) <= '0';
partial_product_25(59) <= '0';
partial_product_25(60) <= '0';
partial_product_25(61) <= '0';
partial_product_25(62) <= '0';
partial_product_25(63) <= '0';
partial_product_25(64) <= '0';
partial_product_25(65) <= '0';
partial_product_25(66) <= '0';
partial_product_25(67) <= '0';
partial_product_25(68) <= '0';
partial_product_25(69) <= '0';
partial_product_25(70) <= '0';
partial_product_25(71) <= '0';
partial_product_25(72) <= '0';
partial_product_25(73) <= '0';
partial_product_25(74) <= '0';
partial_product_25(75) <= '0';
partial_product_25(76) <= '0';
partial_product_25(77) <= '0';
partial_product_25(78) <= '0';
partial_product_25(79) <= '0';
partial_product_25(80) <= '0';
partial_product_25(81) <= '0';
partial_product_25(82) <= '0';
partial_product_25(83) <= '0';
partial_product_25(84) <= '0';
partial_product_25(85) <= '0';
partial_product_25(86) <= '0';
partial_product_25(87) <= '0';
partial_product_25(88) <= '0';
partial_product_25(89) <= '0';
partial_product_25(90) <= '0';
partial_product_25(91) <= '0';
partial_product_25(92) <= '0';
partial_product_25(93) <= '0';
partial_product_25(94) <= '0';
partial_product_25(95) <= '0';
partial_product_25(96) <= '0';
partial_product_25(97) <= '0';
partial_product_25(98) <= '0';
partial_product_25(99) <= '0';
partial_product_25(100) <= '0';
partial_product_25(101) <= '0';
partial_product_25(102) <= '0';
partial_product_25(103) <= '0';
partial_product_25(104) <= '0';
partial_product_25(105) <= '0';
partial_product_25(106) <= '0';
partial_product_25(107) <= '0';
partial_product_25(108) <= '0';
partial_product_25(109) <= '0';
partial_product_25(110) <= '0';
partial_product_25(111) <= '0';
partial_product_25(112) <= '0';
partial_product_25(113) <= '0';
partial_product_25(114) <= '0';
partial_product_25(115) <= '0';
partial_product_25(116) <= '0';
partial_product_25(117) <= '0';
partial_product_25(118) <= '0';
partial_product_25(119) <= '0';
partial_product_25(120) <= '0';
partial_product_25(121) <= '0';
partial_product_25(122) <= '0';
partial_product_25(123) <= '0';
partial_product_25(124) <= '0';
partial_product_25(125) <= '0';
partial_product_25(126) <= '0';
partial_product_25(127) <= '0';
partial_product_25(128) <= '0';
partial_product_25(129) <= '0';
partial_product_25(130) <= '0';
partial_product_25(131) <= '0';
partial_product_25(132) <= '0';
partial_product_25(133) <= '0';
partial_product_25(134) <= '0';
partial_product_25(135) <= '0';
partial_product_25(136) <= '0';
partial_product_25(137) <= '0';
partial_product_25(138) <= '0';
partial_product_25(139) <= '0';
partial_product_25(140) <= '0';
partial_product_25(141) <= '0';
partial_product_25(142) <= '0';
partial_product_25(143) <= '0';
partial_product_25(144) <= '0';
partial_product_25(145) <= '0';
partial_product_25(146) <= '0';
partial_product_25(147) <= '0';
partial_product_25(148) <= '0';
partial_product_25(149) <= '0';
partial_product_25(150) <= '0';
partial_product_25(151) <= '0';
partial_product_25(152) <= '0';
partial_product_25(153) <= '0';
partial_product_25(154) <= '0';
partial_product_25(155) <= '0';
partial_product_25(156) <= '0';
partial_product_25(157) <= '0';
partial_product_25(158) <= '0';
partial_product_25(159) <= '0';
partial_product_25(160) <= '0';
partial_product_25(161) <= '0';
partial_product_25(162) <= '0';
partial_product_25(163) <= '0';
partial_product_25(164) <= '0';
partial_product_25(165) <= '0';
partial_product_25(166) <= '0';
partial_product_25(167) <= '0';
partial_product_25(168) <= '0';
partial_product_25(169) <= '0';
partial_product_25(170) <= '0';
partial_product_25(171) <= '0';
partial_product_25(172) <= '0';
partial_product_25(173) <= '0';
partial_product_25(174) <= '0';
partial_product_25(175) <= '0';
partial_product_25(176) <= '0';
partial_product_25(177) <= '0';
partial_product_25(178) <= '0';
partial_product_25(179) <= '0';
partial_product_25(180) <= '0';
partial_product_25(181) <= '0';
partial_product_25(182) <= '0';
partial_product_25(183) <= '0';
partial_product_25(184) <= '0';
partial_product_25(185) <= '0';
partial_product_25(186) <= '0';
partial_product_25(187) <= '0';
partial_product_25(188) <= '0';
partial_product_25(189) <= '0';
partial_product_25(190) <= '0';
partial_product_25(191) <= '0';
partial_product_25(192) <= '0';
partial_product_25(193) <= '0';
partial_product_25(194) <= '0';
partial_product_25(195) <= '0';
partial_product_25(196) <= '0';
partial_product_25(197) <= '0';
partial_product_25(198) <= '0';
partial_product_25(199) <= '0';
partial_product_25(200) <= '0';
partial_product_25(201) <= '0';
partial_product_25(202) <= '0';
partial_product_25(203) <= '0';
partial_product_25(204) <= '0';
partial_product_25(205) <= '0';
partial_product_25(206) <= '0';
partial_product_25(207) <= '0';
partial_product_25(208) <= '0';
partial_product_25(209) <= '0';
partial_product_25(210) <= '0';
partial_product_25(211) <= '0';
partial_product_25(212) <= '0';
partial_product_25(213) <= '0';
partial_product_25(214) <= '0';
partial_product_25(215) <= '0';
partial_product_25(216) <= '0';
partial_product_25(217) <= '0';
partial_product_25(218) <= '0';
partial_product_25(219) <= '0';
partial_product_25(220) <= '0';
partial_product_25(221) <= '0';
partial_product_25(222) <= '0';
partial_product_25(223) <= '0';
partial_product_25(224) <= '0';
partial_product_25(225) <= '0';
partial_product_25(226) <= '0';
partial_product_25(227) <= '0';
partial_product_25(228) <= '0';
partial_product_25(229) <= '0';
partial_product_25(230) <= '0';
partial_product_25(231) <= '0';
partial_product_25(232) <= '0';
partial_product_25(233) <= '0';
partial_product_25(234) <= '0';
partial_product_25(235) <= '0';
partial_product_25(236) <= '0';
partial_product_25(237) <= '0';
partial_product_25(238) <= '0';
partial_product_25(239) <= '0';
partial_product_25(240) <= '0';
partial_product_25(241) <= '0';
partial_product_25(242) <= '0';
partial_product_25(243) <= '0';
partial_product_25(244) <= '0';
partial_product_25(245) <= '0';
partial_product_25(246) <= '0';
partial_product_25(247) <= '0';
partial_product_25(248) <= '0';
partial_product_25(249) <= '0';
partial_product_25(250) <= '0';
partial_product_25(251) <= '0';
partial_product_25(252) <= '0';
partial_product_25(253) <= '0';
partial_product_25(254) <= '0';
partial_product_25(255) <= temp_mult_87(255);
partial_product_25(256) <= temp_mult_87(256);
partial_product_25(257) <= temp_mult_87(257);
partial_product_25(258) <= temp_mult_87(258);
partial_product_25(259) <= temp_mult_87(259);
partial_product_25(260) <= temp_mult_87(260);
partial_product_25(261) <= temp_mult_87(261);
partial_product_25(262) <= temp_mult_87(262);
partial_product_25(263) <= temp_mult_87(263);
partial_product_25(264) <= temp_mult_87(264);
partial_product_25(265) <= temp_mult_87(265);
partial_product_25(266) <= temp_mult_87(266);
partial_product_25(267) <= temp_mult_87(267);
partial_product_25(268) <= temp_mult_87(268);
partial_product_25(269) <= temp_mult_87(269);
partial_product_25(270) <= temp_mult_87(270);
partial_product_25(271) <= temp_mult_87(271);
partial_product_25(272) <= temp_mult_87(272);
partial_product_25(273) <= temp_mult_87(273);
partial_product_25(274) <= temp_mult_87(274);
partial_product_25(275) <= temp_mult_87(275);
partial_product_25(276) <= temp_mult_87(276);
partial_product_25(277) <= temp_mult_87(277);
partial_product_25(278) <= temp_mult_87(278);
partial_product_25(279) <= temp_mult_87(279);
partial_product_25(280) <= temp_mult_87(280);
partial_product_25(281) <= temp_mult_87(281);
partial_product_25(282) <= temp_mult_87(282);
partial_product_25(283) <= temp_mult_87(283);
partial_product_25(284) <= temp_mult_87(284);
partial_product_25(285) <= temp_mult_87(285);
partial_product_25(286) <= temp_mult_87(286);
partial_product_25(287) <= temp_mult_87(287);
partial_product_25(288) <= temp_mult_87(288);
partial_product_25(289) <= temp_mult_87(289);
partial_product_25(290) <= temp_mult_87(290);
partial_product_25(291) <= temp_mult_87(291);
partial_product_25(292) <= temp_mult_87(292);
partial_product_25(293) <= temp_mult_87(293);
partial_product_25(294) <= temp_mult_87(294);
partial_product_25(295) <= temp_mult_87(295);
partial_product_25(296) <= '0';
partial_product_25(297) <= '0';
partial_product_25(298) <= '0';
partial_product_25(299) <= '0';
partial_product_25(300) <= '0';
partial_product_25(301) <= '0';
partial_product_25(302) <= '0';
partial_product_25(303) <= '0';
partial_product_25(304) <= '0';
partial_product_25(305) <= '0';
partial_product_25(306) <= '0';
partial_product_25(307) <= '0';
partial_product_25(308) <= '0';
partial_product_25(309) <= '0';
partial_product_25(310) <= '0';
partial_product_25(311) <= '0';
partial_product_25(312) <= '0';
partial_product_25(313) <= '0';
partial_product_25(314) <= '0';
partial_product_25(315) <= '0';
partial_product_25(316) <= '0';
partial_product_25(317) <= '0';
partial_product_25(318) <= '0';
partial_product_25(319) <= '0';
partial_product_25(320) <= '0';
partial_product_25(321) <= '0';
partial_product_25(322) <= '0';
partial_product_25(323) <= '0';
partial_product_25(324) <= '0';
partial_product_25(325) <= '0';
partial_product_25(326) <= '0';
partial_product_25(327) <= '0';
partial_product_25(328) <= '0';
partial_product_25(329) <= '0';
partial_product_25(330) <= '0';
partial_product_25(331) <= '0';
partial_product_25(332) <= '0';
partial_product_25(333) <= '0';
partial_product_25(334) <= '0';
partial_product_25(335) <= '0';
partial_product_25(336) <= '0';
partial_product_25(337) <= '0';
partial_product_25(338) <= '0';
partial_product_25(339) <= '0';
partial_product_25(340) <= '0';
partial_product_25(341) <= '0';
partial_product_25(342) <= '0';
partial_product_25(343) <= '0';
partial_product_25(344) <= '0';
partial_product_25(345) <= '0';
partial_product_25(346) <= '0';
partial_product_25(347) <= '0';
partial_product_25(348) <= '0';
partial_product_25(349) <= '0';
partial_product_25(350) <= '0';
partial_product_25(351) <= '0';
partial_product_25(352) <= '0';
partial_product_25(353) <= '0';
partial_product_25(354) <= '0';
partial_product_25(355) <= '0';
partial_product_25(356) <= '0';
partial_product_25(357) <= '0';
partial_product_25(358) <= '0';
partial_product_25(359) <= '0';
partial_product_25(360) <= '0';
partial_product_25(361) <= '0';
partial_product_25(362) <= '0';
partial_product_25(363) <= '0';
partial_product_25(364) <= '0';
partial_product_25(365) <= '0';
partial_product_25(366) <= '0';
partial_product_25(367) <= '0';
partial_product_25(368) <= '0';
partial_product_25(369) <= '0';
partial_product_25(370) <= '0';
partial_product_25(371) <= '0';
partial_product_25(372) <= '0';
partial_product_25(373) <= '0';
partial_product_25(374) <= '0';
partial_product_25(375) <= '0';
partial_product_25(376) <= '0';
partial_product_25(377) <= '0';
partial_product_25(378) <= '0';
partial_product_25(379) <= '0';
partial_product_25(380) <= '0';
partial_product_25(381) <= '0';
partial_product_25(382) <= '0';
partial_product_25(383) <= '0';
partial_product_25(384) <= '0';
partial_product_25(385) <= '0';
partial_product_25(386) <= '0';
partial_product_25(387) <= '0';
partial_product_25(388) <= '0';
partial_product_25(389) <= '0';
partial_product_25(390) <= '0';
partial_product_25(391) <= '0';
partial_product_25(392) <= '0';
partial_product_25(393) <= '0';
partial_product_25(394) <= '0';
partial_product_25(395) <= '0';
partial_product_25(396) <= '0';
partial_product_25(397) <= '0';
partial_product_25(398) <= '0';
partial_product_25(399) <= '0';
partial_product_25(400) <= '0';
partial_product_25(401) <= '0';
partial_product_25(402) <= '0';
partial_product_25(403) <= '0';
partial_product_25(404) <= '0';
partial_product_25(405) <= '0';
partial_product_25(406) <= '0';
partial_product_25(407) <= '0';
partial_product_25(408) <= '0';
partial_product_25(409) <= '0';
partial_product_25(410) <= '0';
partial_product_25(411) <= '0';
partial_product_25(412) <= '0';
partial_product_25(413) <= '0';
partial_product_25(414) <= '0';
partial_product_25(415) <= '0';
partial_product_25(416) <= '0';
partial_product_25(417) <= '0';
partial_product_25(418) <= '0';
partial_product_25(419) <= '0';
partial_product_25(420) <= '0';
partial_product_25(421) <= '0';
partial_product_25(422) <= '0';
partial_product_25(423) <= '0';
partial_product_25(424) <= '0';
partial_product_25(425) <= '0';
partial_product_25(426) <= '0';
partial_product_25(427) <= '0';
partial_product_25(428) <= '0';
partial_product_25(429) <= '0';
partial_product_25(430) <= '0';
partial_product_25(431) <= '0';
partial_product_25(432) <= '0';
partial_product_25(433) <= '0';
partial_product_25(434) <= '0';
partial_product_25(435) <= '0';
partial_product_25(436) <= '0';
partial_product_25(437) <= '0';
partial_product_25(438) <= '0';
partial_product_25(439) <= '0';
partial_product_25(440) <= '0';
partial_product_25(441) <= '0';
partial_product_25(442) <= '0';
partial_product_25(443) <= '0';
partial_product_25(444) <= '0';
partial_product_25(445) <= '0';
partial_product_25(446) <= '0';
partial_product_25(447) <= '0';
partial_product_25(448) <= '0';
partial_product_25(449) <= '0';
partial_product_25(450) <= '0';
partial_product_25(451) <= '0';
partial_product_25(452) <= '0';
partial_product_25(453) <= '0';
partial_product_25(454) <= '0';
partial_product_25(455) <= '0';
partial_product_25(456) <= '0';
partial_product_25(457) <= '0';
partial_product_25(458) <= '0';
partial_product_25(459) <= '0';
partial_product_25(460) <= '0';
partial_product_25(461) <= '0';
partial_product_25(462) <= '0';
partial_product_25(463) <= '0';
partial_product_25(464) <= '0';
partial_product_25(465) <= '0';
partial_product_25(466) <= '0';
partial_product_25(467) <= '0';
partial_product_25(468) <= '0';
partial_product_25(469) <= '0';
partial_product_25(470) <= '0';
partial_product_25(471) <= '0';
partial_product_25(472) <= '0';
partial_product_25(473) <= '0';
partial_product_25(474) <= '0';
partial_product_25(475) <= '0';
partial_product_25(476) <= '0';
partial_product_25(477) <= '0';
partial_product_25(478) <= '0';
partial_product_25(479) <= '0';
partial_product_25(480) <= '0';
partial_product_25(481) <= '0';
partial_product_25(482) <= '0';
partial_product_25(483) <= '0';
partial_product_25(484) <= '0';
partial_product_25(485) <= '0';
partial_product_25(486) <= '0';
partial_product_25(487) <= '0';
partial_product_25(488) <= '0';
partial_product_25(489) <= '0';
partial_product_25(490) <= '0';
partial_product_25(491) <= '0';
partial_product_25(492) <= '0';
partial_product_25(493) <= '0';
partial_product_25(494) <= '0';
partial_product_25(495) <= '0';
partial_product_25(496) <= '0';
partial_product_25(497) <= '0';
partial_product_25(498) <= '0';
partial_product_25(499) <= '0';
partial_product_25(500) <= '0';
partial_product_25(501) <= '0';
partial_product_25(502) <= '0';
partial_product_25(503) <= '0';
partial_product_25(504) <= '0';
partial_product_25(505) <= '0';
partial_product_25(506) <= '0';
partial_product_25(507) <= '0';
partial_product_25(508) <= '0';
partial_product_25(509) <= '0';
partial_product_25(510) <= '0';
partial_product_25(511) <= '0';
partial_product_25(512) <= '0';

partial_product_26(255 downto 0) <= (others => '0');
partial_product_26(513 downto 256) <= temp_mult_161;

partial_product_27(255 downto 0) <= (others => '0');
partial_product_27(513 downto 256) <= temp_mult_162;

process(clk)
begin
    if(rising_edge(clk)) then
        temp_comp_1_a1  <= "0" & partial_product_0;
        temp_comp_1_a2  <= "0" & partial_product_1;
        temp_comp_1_a3  <= "0" & partial_product_2;
        temp_comp_1_a4  <= "0" & partial_product_3;
        temp_comp_1_a5  <= "0" & partial_product_4;
        temp_comp_1_a6  <= "0" & partial_product_5;
        temp_comp_1_a7  <= "0" & partial_product_6;
        temp_comp_1_a8  <= "0" & partial_product_7;
        temp_comp_1_a9  <= "0" & partial_product_8;
        temp_comp_1_a10 <= "0" & partial_product_9;
        temp_comp_1_a11 <= "0" & partial_product_10;
        temp_comp_1_a12 <= "0" & partial_product_11;
        temp_comp_1_a13 <= "0" & partial_product_12;
        temp_comp_1_a14 <= "0" & partial_product_13;
        temp_comp_1_a15 <= "0" & partial_product_14;
        temp_comp_1_a16 <= "0" & partial_product_15;
        temp_comp_1_a17 <= "0" & partial_product_16;
        temp_comp_1_a18 <= "0" & partial_product_17;
        temp_comp_1_a19 <= "0" & partial_product_18;
        temp_comp_1_a20 <= "0" & partial_product_19;
        temp_comp_1_a21 <= "0" & partial_product_20;
        temp_comp_1_a22 <= "0" & partial_product_21;
        temp_comp_1_a23 <= "0" & partial_product_22;
        temp_comp_1_a24 <= "0" & partial_product_23;
        temp_comp_1_a25 <= "0" & partial_product_24;
        temp_comp_1_a26 <= "0" & partial_product_25;
        temp_comp_1_a27 <= not partial_product_26;
        temp_comp_1_a28 <= not partial_product_27;
        temp_comp_1_a29(0) <= '1';
        temp_comp_1_a29(513 downto 1) <= (others => '0');
        temp_comp_1_a30(0) <= '1';
        temp_comp_1_a30(513 downto 1) <= (others => '0');
    end if;
end process;

temp_comp_1 : adder_compressor_30_5
    Generic Map(
        total_size => 514
    )
    Port Map(
        a1 => temp_comp_1_a1,
        a2 => temp_comp_1_a2,
        a3 => temp_comp_1_a3,
        a4 => temp_comp_1_a4,
        a5 => temp_comp_1_a5,
        a6 => temp_comp_1_a6,
        a7 => temp_comp_1_a7,
        a8 => temp_comp_1_a8,
        a9 => temp_comp_1_a9,
        a10=> temp_comp_1_a10,
        a11=> temp_comp_1_a11,
        a12=> temp_comp_1_a12,
        a13=> temp_comp_1_a13,
        a14=> temp_comp_1_a14,
        a15=> temp_comp_1_a15,
        a16=> temp_comp_1_a16,
        a17=> temp_comp_1_a17,
        a18=> temp_comp_1_a18,
        a19=> temp_comp_1_a19,
        a20=> temp_comp_1_a20,
        a21=> temp_comp_1_a21,
        a22=> temp_comp_1_a22,
        a23=> temp_comp_1_a23,
        a24=> temp_comp_1_a24,
        a25=> temp_comp_1_a25,
        a26=> temp_comp_1_a26,
        a27=> temp_comp_1_a27,
        a28=> temp_comp_1_a28,
        a29=> temp_comp_1_a29,
        a30=> temp_comp_1_a30,
        c1 => temp_comp_1_c1,
        c2 => temp_comp_1_c2,
        c3 => temp_comp_1_c3,
        c4 => temp_comp_1_c4,
        s  => temp_comp_1_s
    );

process(clk)
begin
    if(rising_edge(clk)) then
        temp_comp_2_a1 <= temp_comp_1_c1(513 downto 0);
        temp_comp_2_a2 <= temp_comp_1_c2(513 downto 0);
        temp_comp_2_a3 <= temp_comp_1_c3(513 downto 0);
        temp_comp_2_a4 <= temp_comp_1_c4(513 downto 0);
        temp_comp_2_a5 <= temp_comp_1_s(513 downto 0);
    end if;
end process;

temp_comp_2 : adder_compressor_5_3
    Generic Map(
        total_size => 514
    )
    Port Map(
        a1 => temp_comp_2_a1,
        a2 => temp_comp_2_a2,
        a3 => temp_comp_2_a3,
        a4 => temp_comp_2_a4,
        a5 => temp_comp_2_a5,
        c1 => temp_comp_2_c1,
        c2 => temp_comp_2_c2,
        s => temp_comp_2_s
    );

temp_comp_3_a1 <= temp_comp_2_c1(513 downto 0);
temp_comp_3_a2 <= temp_comp_2_c2(513 downto 0);
temp_comp_3_a3 <= temp_comp_2_s(513 downto 0);

temp_comp_3 : adder_compressor_3_2
    Generic Map(
        total_size => 514
    )
    Port Map(
        a => temp_comp_3_a1,
        b => temp_comp_3_a2,
        p => temp_comp_3_a3,
        c => temp_comp_3_c,
        s => temp_comp_3_s
    );

process(clk)
begin
    if(rising_edge(clk)) then
        temp_comp_4_a1 <= temp_comp_3_c(513 downto 0);
        temp_comp_4_a2 <= temp_comp_3_s(513 downto 0);
    end if;
end process;

final_comp_a <= temp_comp_4_a1;
final_comp_b <= temp_comp_4_a2;

final_comp : entity work.wide_adder_carry_select(behavioral_aam)
    Generic Map(
        base_size => 2,
        total_size => 514
    )
    Port Map(
        a => final_comp_a,
        b => final_comp_b,
        cin => "0",
        o => final_comp_o
    );

process(clk)
begin
    if(rising_edge(clk)) then
        temp_o4 <= unsigned(final_comp_o);
        o <= std_logic_vector(temp_o4);
    end if;
end process;

end tiled_behavioral_v2;